magic
tech sky130A
magscale 1 2
timestamp 1672276304
<< viali >>
rect 3617 57545 3651 57579
rect 5641 57545 5675 57579
rect 10333 57545 10367 57579
rect 11713 57545 11747 57579
rect 13093 57545 13127 57579
rect 14473 57545 14507 57579
rect 15853 57545 15887 57579
rect 17233 57545 17267 57579
rect 18613 57545 18647 57579
rect 19993 57545 20027 57579
rect 21373 57545 21407 57579
rect 22753 57545 22787 57579
rect 29101 57545 29135 57579
rect 29837 57545 29871 57579
rect 30573 57545 30607 57579
rect 40049 57545 40083 57579
rect 42165 57545 42199 57579
rect 51273 57545 51307 57579
rect 4261 57477 4295 57511
rect 45845 57477 45879 57511
rect 52653 57477 52687 57511
rect 5825 57409 5859 57443
rect 6377 57409 6411 57443
rect 7481 57409 7515 57443
rect 8309 57409 8343 57443
rect 9137 57409 9171 57443
rect 10517 57409 10551 57443
rect 11897 57409 11931 57443
rect 13277 57409 13311 57443
rect 14657 57409 14691 57443
rect 16037 57409 16071 57443
rect 17417 57409 17451 57443
rect 18797 57409 18831 57443
rect 20177 57409 20211 57443
rect 21557 57409 21591 57443
rect 22937 57409 22971 57443
rect 24133 57409 24167 57443
rect 24317 57409 24351 57443
rect 25329 57409 25363 57443
rect 25513 57409 25547 57443
rect 26893 57409 26927 57443
rect 27905 57409 27939 57443
rect 29285 57409 29319 57443
rect 30389 57409 30423 57443
rect 31769 57409 31803 57443
rect 33333 57409 33367 57443
rect 34529 57409 34563 57443
rect 34713 57409 34747 57443
rect 34989 57409 35023 57443
rect 36185 57409 36219 57443
rect 37565 57409 37599 57443
rect 38669 57409 38703 57443
rect 40417 57409 40451 57443
rect 41981 57409 42015 57443
rect 42257 57409 42291 57443
rect 44373 57409 44407 57443
rect 46949 57409 46983 57443
rect 48329 57409 48363 57443
rect 48605 57409 48639 57443
rect 49709 57409 49743 57443
rect 51457 57409 51491 57443
rect 53941 57409 53975 57443
rect 55321 57409 55355 57443
rect 56609 57409 56643 57443
rect 23949 57341 23983 57375
rect 26709 57341 26743 57375
rect 27629 57341 27663 57375
rect 32045 57341 32079 57375
rect 33609 57341 33643 57375
rect 35909 57341 35943 57375
rect 37289 57341 37323 57375
rect 38945 57341 38979 57375
rect 40233 57341 40267 57375
rect 40325 57341 40359 57375
rect 40509 57341 40543 57375
rect 42809 57341 42843 57375
rect 43085 57341 43119 57375
rect 44649 57341 44683 57375
rect 47225 57341 47259 57375
rect 49985 57341 50019 57375
rect 4445 57273 4479 57307
rect 27813 57273 27847 57307
rect 33149 57273 33183 57307
rect 33517 57273 33551 57307
rect 55505 57273 55539 57307
rect 11161 57205 11195 57239
rect 20821 57205 20855 57239
rect 22109 57205 22143 57239
rect 25697 57205 25731 57239
rect 27077 57205 27111 57239
rect 27721 57205 27755 57239
rect 28457 57205 28491 57239
rect 31125 57205 31159 57239
rect 34897 57205 34931 57239
rect 41797 57205 41831 57239
rect 44189 57205 44223 57239
rect 44557 57205 44591 57239
rect 45753 57205 45787 57239
rect 52745 57205 52779 57239
rect 54125 57205 54159 57239
rect 4721 57001 4755 57035
rect 5917 57001 5951 57035
rect 6561 57001 6595 57035
rect 8861 57001 8895 57035
rect 10241 57001 10275 57035
rect 11621 57001 11655 57035
rect 13001 57001 13035 57035
rect 14381 57001 14415 57035
rect 15761 57001 15795 57035
rect 17141 57001 17175 57035
rect 18521 57001 18555 57035
rect 19901 57001 19935 57035
rect 21281 57001 21315 57035
rect 23029 57001 23063 57035
rect 24317 57001 24351 57035
rect 27077 57001 27111 57035
rect 28089 57001 28123 57035
rect 34253 57001 34287 57035
rect 37289 57001 37323 57035
rect 47593 57001 47627 57035
rect 48881 57001 48915 57035
rect 49709 57001 49743 57035
rect 50353 57001 50387 57035
rect 50997 57001 51031 57035
rect 51641 57001 51675 57035
rect 52469 57001 52503 57035
rect 53113 57001 53147 57035
rect 53757 57001 53791 57035
rect 54401 57001 54435 57035
rect 56241 57001 56275 57035
rect 22293 56933 22327 56967
rect 27629 56933 27663 56967
rect 42901 56933 42935 56967
rect 44281 56933 44315 56967
rect 48237 56933 48271 56967
rect 23673 56865 23707 56899
rect 25697 56865 25731 56899
rect 26433 56865 26467 56899
rect 26525 56865 26559 56899
rect 31125 56865 31159 56899
rect 35173 56865 35207 56899
rect 36185 56865 36219 56899
rect 38669 56865 38703 56899
rect 39037 56865 39071 56899
rect 39129 56865 39163 56899
rect 40785 56865 40819 56899
rect 42993 56865 43027 56899
rect 44189 56865 44223 56899
rect 45017 56865 45051 56899
rect 55229 56865 55263 56899
rect 22477 56797 22511 56831
rect 23213 56797 23247 56831
rect 23765 56797 23799 56831
rect 24192 56797 24226 56831
rect 25326 56797 25360 56831
rect 25789 56797 25823 56831
rect 26952 56797 26986 56831
rect 27813 56797 27847 56831
rect 27905 56797 27939 56831
rect 28181 56797 28215 56831
rect 29285 56797 29319 56831
rect 29469 56797 29503 56831
rect 29561 56797 29595 56831
rect 29653 56797 29687 56831
rect 29837 56797 29871 56831
rect 30941 56797 30975 56831
rect 31033 56797 31067 56831
rect 31217 56797 31251 56831
rect 31950 56797 31984 56831
rect 32321 56797 32355 56831
rect 32413 56797 32447 56831
rect 33425 56797 33459 56831
rect 33517 56797 33551 56831
rect 33701 56797 33735 56831
rect 33793 56797 33827 56831
rect 34437 56797 34471 56831
rect 34621 56797 34655 56831
rect 34713 56797 34747 56831
rect 36001 56797 36035 56831
rect 36553 56797 36587 56831
rect 36829 56797 36863 56831
rect 37473 56797 37507 56831
rect 37749 56797 37783 56831
rect 38853 56797 38887 56831
rect 38945 56797 38979 56831
rect 39773 56797 39807 56831
rect 40358 56797 40392 56831
rect 40877 56797 40911 56831
rect 41705 56797 41739 56831
rect 41797 56797 41831 56831
rect 41981 56797 42015 56831
rect 42073 56797 42107 56831
rect 42533 56797 42567 56831
rect 42717 56797 42751 56831
rect 43453 56797 43487 56831
rect 44373 56797 44407 56831
rect 44741 56797 44775 56831
rect 45661 56797 45695 56831
rect 46121 56797 46155 56831
rect 46949 56797 46983 56831
rect 24133 56661 24167 56695
rect 25145 56661 25179 56695
rect 25329 56661 25363 56695
rect 26893 56661 26927 56695
rect 29101 56661 29135 56695
rect 30757 56661 30791 56695
rect 31769 56661 31803 56695
rect 31953 56661 31987 56695
rect 33241 56661 33275 56695
rect 36093 56661 36127 56695
rect 37657 56661 37691 56695
rect 40233 56661 40267 56695
rect 40417 56661 40451 56695
rect 41521 56661 41555 56695
rect 45477 56661 45511 56695
rect 24041 56457 24075 56491
rect 28089 56457 28123 56491
rect 31769 56457 31803 56491
rect 32689 56457 32723 56491
rect 35541 56457 35575 56491
rect 36369 56457 36403 56491
rect 37289 56457 37323 56491
rect 49249 56457 49283 56491
rect 51089 56457 51123 56491
rect 51641 56457 51675 56491
rect 52469 56457 52503 56491
rect 53849 56457 53883 56491
rect 55229 56457 55263 56491
rect 28457 56389 28491 56423
rect 33885 56389 33919 56423
rect 34713 56389 34747 56423
rect 36737 56389 36771 56423
rect 40417 56389 40451 56423
rect 22661 56321 22695 56355
rect 24225 56321 24259 56355
rect 25513 56321 25547 56355
rect 26259 56321 26293 56355
rect 27353 56321 27387 56355
rect 28273 56321 28307 56355
rect 29193 56321 29227 56355
rect 29377 56321 29411 56355
rect 29469 56321 29503 56355
rect 29653 56321 29687 56355
rect 30297 56321 30331 56355
rect 30941 56321 30975 56355
rect 31953 56321 31987 56355
rect 32229 56321 32263 56355
rect 32873 56321 32907 56355
rect 34529 56321 34563 56355
rect 34805 56321 34839 56355
rect 35265 56321 35299 56355
rect 35633 56321 35667 56355
rect 35725 56321 35759 56355
rect 36553 56321 36587 56355
rect 37657 56321 37691 56355
rect 39221 56321 39255 56355
rect 39313 56321 39347 56355
rect 39497 56321 39531 56355
rect 40187 56321 40221 56355
rect 40325 56321 40359 56355
rect 40509 56321 40543 56355
rect 41397 56321 41431 56355
rect 41521 56321 41555 56355
rect 42165 56321 42199 56355
rect 42257 56321 42291 56355
rect 43177 56321 43211 56355
rect 44005 56321 44039 56355
rect 44281 56321 44315 56355
rect 44833 56321 44867 56355
rect 46857 56321 46891 56355
rect 47501 56321 47535 56355
rect 48329 56321 48363 56355
rect 23581 56253 23615 56287
rect 24409 56253 24443 56287
rect 25329 56253 25363 56287
rect 26525 56253 26559 56287
rect 27537 56253 27571 56287
rect 30481 56253 30515 56287
rect 33149 56253 33183 56287
rect 37749 56253 37783 56287
rect 38301 56253 38335 56287
rect 38761 56253 38795 56287
rect 40049 56253 40083 56287
rect 41613 56253 41647 56287
rect 43085 56253 43119 56287
rect 43821 56253 43855 56287
rect 45569 56253 45603 56287
rect 29285 56185 29319 56219
rect 38393 56185 38427 56219
rect 40693 56185 40727 56219
rect 42809 56185 42843 56219
rect 44097 56185 44131 56219
rect 44189 56185 44223 56219
rect 46213 56185 46247 56219
rect 25697 56117 25731 56151
rect 27169 56117 27203 56151
rect 29009 56117 29043 56151
rect 30113 56117 30147 56151
rect 32137 56117 32171 56151
rect 33057 56117 33091 56151
rect 33793 56117 33827 56151
rect 34529 56117 34563 56151
rect 39497 56117 39531 56151
rect 41153 56117 41187 56151
rect 23121 55913 23155 55947
rect 23673 55913 23707 55947
rect 24133 55913 24167 55947
rect 26065 55913 26099 55947
rect 34253 55913 34287 55947
rect 35265 55913 35299 55947
rect 39221 55913 39255 55947
rect 40509 55913 40543 55947
rect 43637 55913 43671 55947
rect 44373 55913 44407 55947
rect 45661 55913 45695 55947
rect 46949 55913 46983 55947
rect 47869 55913 47903 55947
rect 27077 55845 27111 55879
rect 28641 55845 28675 55879
rect 40141 55845 40175 55879
rect 29009 55777 29043 55811
rect 29101 55777 29135 55811
rect 33517 55777 33551 55811
rect 34621 55777 34655 55811
rect 36829 55777 36863 55811
rect 37197 55777 37231 55811
rect 40049 55777 40083 55811
rect 46397 55777 46431 55811
rect 24317 55709 24351 55743
rect 25237 55709 25271 55743
rect 25881 55709 25915 55743
rect 26801 55709 26835 55743
rect 28825 55709 28859 55743
rect 28917 55709 28951 55743
rect 29653 55709 29687 55743
rect 30849 55709 30883 55743
rect 31125 55709 31159 55743
rect 31309 55709 31343 55743
rect 32137 55709 32171 55743
rect 32413 55709 32447 55743
rect 33149 55709 33183 55743
rect 33333 55709 33367 55743
rect 34451 55709 34485 55743
rect 35357 55709 35391 55743
rect 36184 55709 36218 55743
rect 36277 55709 36311 55743
rect 37013 55709 37047 55743
rect 37657 55709 37691 55743
rect 37841 55709 37875 55743
rect 38117 55709 38151 55743
rect 38669 55709 38703 55743
rect 38775 55709 38809 55743
rect 38945 55709 38979 55743
rect 39037 55709 39071 55743
rect 40325 55709 40359 55743
rect 41613 55709 41647 55743
rect 41889 55709 41923 55743
rect 42533 55709 42567 55743
rect 42625 55687 42659 55721
rect 42753 55709 42787 55743
rect 44464 55709 44498 55743
rect 44557 55709 44591 55743
rect 45201 55709 45235 55743
rect 27077 55641 27111 55675
rect 27997 55641 28031 55675
rect 28181 55641 28215 55675
rect 30987 55641 31021 55675
rect 31217 55641 31251 55675
rect 31953 55641 31987 55675
rect 43269 55641 43303 55675
rect 43453 55641 43487 55675
rect 25421 55573 25455 55607
rect 26893 55573 26927 55607
rect 27813 55573 27847 55607
rect 29837 55573 29871 55607
rect 31493 55573 31527 55607
rect 32321 55573 32355 55607
rect 35909 55573 35943 55607
rect 38025 55573 38059 55607
rect 41429 55573 41463 55607
rect 41797 55573 41831 55607
rect 42349 55573 42383 55607
rect 45017 55573 45051 55607
rect 25513 55369 25547 55403
rect 30290 55369 30324 55403
rect 30849 55369 30883 55403
rect 34529 55369 34563 55403
rect 38025 55369 38059 55403
rect 41613 55369 41647 55403
rect 44741 55369 44775 55403
rect 45569 55369 45603 55403
rect 46121 55369 46155 55403
rect 27997 55301 28031 55335
rect 30205 55301 30239 55335
rect 31033 55301 31067 55335
rect 25697 55233 25731 55267
rect 27077 55233 27111 55267
rect 29285 55233 29319 55267
rect 29377 55233 29411 55267
rect 29520 55233 29554 55267
rect 29663 55233 29697 55267
rect 30113 55233 30147 55267
rect 30389 55233 30423 55267
rect 31217 55233 31251 55267
rect 31861 55233 31895 55267
rect 33241 55233 33275 55267
rect 34713 55233 34747 55267
rect 34989 55233 35023 55267
rect 38209 55233 38243 55267
rect 39037 55233 39071 55267
rect 40233 55233 40267 55267
rect 42073 55233 42107 55267
rect 43177 55233 43211 55267
rect 44005 55233 44039 55267
rect 44189 55233 44223 55267
rect 44925 55233 44959 55267
rect 24041 55165 24075 55199
rect 25053 55165 25087 55199
rect 26617 55165 26651 55199
rect 29101 55165 29135 55199
rect 33701 55165 33735 55199
rect 35541 55165 35575 55199
rect 38393 55165 38427 55199
rect 39129 55165 39163 55199
rect 41981 55165 42015 55199
rect 43269 55165 43303 55199
rect 43821 55165 43855 55199
rect 44281 55165 44315 55199
rect 27261 55097 27295 55131
rect 28273 55097 28307 55131
rect 34805 55097 34839 55131
rect 34897 55097 34931 55131
rect 36185 55097 36219 55131
rect 37289 55097 37323 55131
rect 42809 55097 42843 55131
rect 28457 55029 28491 55063
rect 31953 55029 31987 55063
rect 32321 55029 32355 55063
rect 32781 55029 32815 55063
rect 33149 55029 33183 55063
rect 39405 55029 39439 55063
rect 40509 55029 40543 55063
rect 40693 55029 40727 55063
rect 42257 55029 42291 55063
rect 25145 54825 25179 54859
rect 25789 54825 25823 54859
rect 26341 54825 26375 54859
rect 26893 54825 26927 54859
rect 28181 54825 28215 54859
rect 29837 54825 29871 54859
rect 30389 54825 30423 54859
rect 31401 54825 31435 54859
rect 34805 54825 34839 54859
rect 36001 54825 36035 54859
rect 36829 54825 36863 54859
rect 38117 54825 38151 54859
rect 38669 54825 38703 54859
rect 39865 54825 39899 54859
rect 41521 54825 41555 54859
rect 43453 54825 43487 54859
rect 44557 54825 44591 54859
rect 29193 54757 29227 54791
rect 32597 54757 32631 54791
rect 42993 54757 43027 54791
rect 28733 54689 28767 54723
rect 30849 54689 30883 54723
rect 32321 54689 32355 54723
rect 33885 54689 33919 54723
rect 34253 54689 34287 54723
rect 35173 54689 35207 54723
rect 36369 54689 36403 54723
rect 40325 54689 40359 54723
rect 41705 54689 41739 54723
rect 25605 54621 25639 54655
rect 27077 54621 27111 54655
rect 27997 54621 28031 54655
rect 28181 54621 28215 54655
rect 28825 54621 28859 54655
rect 30757 54621 30791 54655
rect 32229 54621 32263 54655
rect 33793 54621 33827 54655
rect 35081 54621 35115 54655
rect 35909 54621 35943 54655
rect 36185 54621 36219 54655
rect 37749 54621 37783 54655
rect 37933 54621 37967 54655
rect 38853 54621 38887 54655
rect 39037 54621 39071 54655
rect 39497 54621 39531 54655
rect 39681 54621 39715 54655
rect 40509 54621 40543 54655
rect 40785 54621 40819 54655
rect 41797 54621 41831 54655
rect 42717 54621 42751 54655
rect 42993 54621 43027 54655
rect 40693 54553 40727 54587
rect 42809 54553 42843 54587
rect 33609 54485 33643 54519
rect 26249 54281 26283 54315
rect 29193 54281 29227 54315
rect 30021 54281 30055 54315
rect 31953 54281 31987 54315
rect 32321 54281 32355 54315
rect 32873 54281 32907 54315
rect 33793 54281 33827 54315
rect 36093 54281 36127 54315
rect 36645 54281 36679 54315
rect 40233 54281 40267 54315
rect 41337 54281 41371 54315
rect 41965 54281 41999 54315
rect 43729 54281 43763 54315
rect 30941 54213 30975 54247
rect 33241 54213 33275 54247
rect 34529 54213 34563 54247
rect 40049 54213 40083 54247
rect 42165 54213 42199 54247
rect 26801 54145 26835 54179
rect 28273 54145 28307 54179
rect 29377 54145 29411 54179
rect 29561 54145 29595 54179
rect 30205 54145 30239 54179
rect 30389 54145 30423 54179
rect 30849 54145 30883 54179
rect 31033 54145 31067 54179
rect 32137 54145 32171 54179
rect 32413 54145 32447 54179
rect 33057 54145 33091 54179
rect 33333 54145 33367 54179
rect 33977 54145 34011 54179
rect 34713 54145 34747 54179
rect 34805 54145 34839 54179
rect 34897 54145 34931 54179
rect 35449 54145 35483 54179
rect 37289 54145 37323 54179
rect 37933 54145 37967 54179
rect 38577 54145 38611 54179
rect 39497 54145 39531 54179
rect 40325 54145 40359 54179
rect 40877 54145 40911 54179
rect 42901 54145 42935 54179
rect 28457 54009 28491 54043
rect 40049 54009 40083 54043
rect 27721 53941 27755 53975
rect 40969 53941 41003 53975
rect 41797 53941 41831 53975
rect 41981 53941 42015 53975
rect 28089 53737 28123 53771
rect 28641 53737 28675 53771
rect 29653 53737 29687 53771
rect 30389 53737 30423 53771
rect 31125 53737 31159 53771
rect 31953 53737 31987 53771
rect 33333 53737 33367 53771
rect 33977 53737 34011 53771
rect 35081 53737 35115 53771
rect 36001 53737 36035 53771
rect 37013 53737 37047 53771
rect 38669 53737 38703 53771
rect 39405 53737 39439 53771
rect 40417 53737 40451 53771
rect 41429 53737 41463 53771
rect 41981 53737 42015 53771
rect 33149 53669 33183 53703
rect 37565 53669 37599 53703
rect 39865 53669 39899 53703
rect 32597 53601 32631 53635
rect 34621 53601 34655 53635
rect 36461 53601 36495 53635
rect 29377 53533 29411 53567
rect 29653 53533 29687 53567
rect 33317 53465 33351 53499
rect 33517 53465 33551 53499
rect 29469 53397 29503 53431
rect 29377 53193 29411 53227
rect 30021 53193 30055 53227
rect 30481 53193 30515 53227
rect 32597 53193 32631 53227
rect 33333 53193 33367 53227
rect 40693 53193 40727 53227
rect 34713 53125 34747 53159
rect 33977 52989 34011 53023
rect 34529 52989 34563 53023
rect 34989 52989 35023 53023
rect 35173 52649 35207 52683
rect 30665 8041 30699 8075
rect 31585 8041 31619 8075
rect 29561 7837 29595 7871
rect 29469 7701 29503 7735
rect 27353 7361 27387 7395
rect 29653 7361 29687 7395
rect 30297 7361 30331 7395
rect 30757 7361 30791 7395
rect 32045 7361 32079 7395
rect 32689 7361 32723 7395
rect 27445 7157 27479 7191
rect 27997 7157 28031 7191
rect 29561 7157 29595 7191
rect 30205 7157 30239 7191
rect 30849 7157 30883 7191
rect 32137 7157 32171 7191
rect 32781 7157 32815 7191
rect 31125 6817 31159 6851
rect 25605 6749 25639 6783
rect 26249 6749 26283 6783
rect 26893 6749 26927 6783
rect 27629 6749 27663 6783
rect 28457 6749 28491 6783
rect 29101 6749 29135 6783
rect 29561 6749 29595 6783
rect 30849 6749 30883 6783
rect 31769 6749 31803 6783
rect 32413 6749 32447 6783
rect 33149 6749 33183 6783
rect 33977 6749 34011 6783
rect 25145 6613 25179 6647
rect 26341 6613 26375 6647
rect 32505 6613 32539 6647
rect 25053 6409 25087 6443
rect 26801 6341 26835 6375
rect 29469 6341 29503 6375
rect 32045 6341 32079 6375
rect 25697 6273 25731 6307
rect 29285 6273 29319 6307
rect 31769 6273 31803 6307
rect 34529 6273 34563 6307
rect 26617 6205 26651 6239
rect 27537 6205 27571 6239
rect 30021 6205 30055 6239
rect 32873 6137 32907 6171
rect 25605 6069 25639 6103
rect 33333 6069 33367 6103
rect 34621 6069 34655 6103
rect 26709 5729 26743 5763
rect 28641 5729 28675 5763
rect 30757 5729 30791 5763
rect 30941 5729 30975 5763
rect 31677 5729 31711 5763
rect 33333 5729 33367 5763
rect 34805 5729 34839 5763
rect 34989 5729 35023 5763
rect 23489 5661 23523 5695
rect 24317 5661 24351 5695
rect 25237 5661 25271 5695
rect 27905 5661 27939 5695
rect 25421 5593 25455 5627
rect 28089 5593 28123 5627
rect 24225 5525 24259 5559
rect 25421 5253 25455 5287
rect 26801 5253 26835 5287
rect 29561 5253 29595 5287
rect 33425 5253 33459 5287
rect 36185 5253 36219 5287
rect 24593 5185 24627 5219
rect 25697 5185 25731 5219
rect 26617 5185 26651 5219
rect 29377 5185 29411 5219
rect 33609 5185 33643 5219
rect 24133 5117 24167 5151
rect 27721 5117 27755 5151
rect 30389 5117 30423 5151
rect 31769 5117 31803 5151
rect 34529 5117 34563 5151
rect 36369 5117 36403 5151
rect 22661 4981 22695 5015
rect 24685 4981 24719 5015
rect 37197 4777 37231 4811
rect 22385 4709 22419 4743
rect 23673 4641 23707 4675
rect 25237 4641 25271 4675
rect 25421 4641 25455 4675
rect 26249 4641 26283 4675
rect 27629 4641 27663 4675
rect 27813 4641 27847 4675
rect 28181 4641 28215 4675
rect 30849 4641 30883 4675
rect 33149 4641 33183 4675
rect 33333 4641 33367 4675
rect 33609 4641 33643 4675
rect 20729 4573 20763 4607
rect 21557 4573 21591 4607
rect 23029 4573 23063 4607
rect 24133 4573 24167 4607
rect 30389 4573 30423 4607
rect 36093 4573 36127 4607
rect 36737 4573 36771 4607
rect 37841 4573 37875 4607
rect 30573 4505 30607 4539
rect 22937 4437 22971 4471
rect 24225 4437 24259 4471
rect 36645 4437 36679 4471
rect 36185 4165 36219 4199
rect 22753 4097 22787 4131
rect 26617 4097 26651 4131
rect 29193 4097 29227 4131
rect 32137 4097 32171 4131
rect 36369 4097 36403 4131
rect 21005 4029 21039 4063
rect 23857 4029 23891 4063
rect 24041 4029 24075 4063
rect 25697 4029 25731 4063
rect 26801 4029 26835 4063
rect 28457 4029 28491 4063
rect 29377 4029 29411 4063
rect 29745 4029 29779 4063
rect 32321 4029 32355 4063
rect 32781 4029 32815 4063
rect 34529 4029 34563 4063
rect 37933 4029 37967 4063
rect 40049 4029 40083 4063
rect 21649 3961 21683 3995
rect 38577 3961 38611 3995
rect 40693 3961 40727 3995
rect 17233 3893 17267 3927
rect 18521 3893 18555 3927
rect 19533 3893 19567 3927
rect 20177 3893 20211 3927
rect 22293 3893 22327 3927
rect 22845 3893 22879 3927
rect 37289 3893 37323 3927
rect 39221 3893 39255 3927
rect 20269 3621 20303 3655
rect 38669 3621 38703 3655
rect 41429 3621 41463 3655
rect 43361 3621 43395 3655
rect 19625 3553 19659 3587
rect 22477 3553 22511 3587
rect 22661 3553 22695 3587
rect 25237 3553 25271 3587
rect 27997 3553 28031 3587
rect 28181 3553 28215 3587
rect 28457 3553 28491 3587
rect 31033 3553 31067 3587
rect 33609 3553 33643 3587
rect 36369 3553 36403 3587
rect 39957 3553 39991 3587
rect 42073 3553 42107 3587
rect 10333 3485 10367 3519
rect 12265 3485 12299 3519
rect 13093 3485 13127 3519
rect 14197 3485 14231 3519
rect 15025 3485 15059 3519
rect 15853 3485 15887 3519
rect 16681 3485 16715 3519
rect 17509 3485 17543 3519
rect 18153 3485 18187 3519
rect 18797 3485 18831 3519
rect 20913 3485 20947 3519
rect 21557 3485 21591 3519
rect 30573 3485 30607 3519
rect 33149 3485 33183 3519
rect 35909 3485 35943 3519
rect 39313 3485 39347 3519
rect 40601 3485 40635 3519
rect 42717 3485 42751 3519
rect 44189 3485 44223 3519
rect 45017 3485 45051 3519
rect 46949 3485 46983 3519
rect 47777 3485 47811 3519
rect 49709 3485 49743 3519
rect 50537 3485 50571 3519
rect 52469 3485 52503 3519
rect 24317 3417 24351 3451
rect 25421 3417 25455 3451
rect 27077 3417 27111 3451
rect 30757 3417 30791 3451
rect 33333 3417 33367 3451
rect 36093 3417 36127 3451
rect 22201 3145 22235 3179
rect 24041 3077 24075 3111
rect 25697 3077 25731 3111
rect 21649 3009 21683 3043
rect 22109 3009 22143 3043
rect 23857 3009 23891 3043
rect 37289 3009 37323 3043
rect 41337 3009 41371 3043
rect 17417 2941 17451 2975
rect 20177 2941 20211 2975
rect 21005 2941 21039 2975
rect 26617 2941 26651 2975
rect 26801 2941 26835 2975
rect 28457 2941 28491 2975
rect 29377 2941 29411 2975
rect 29561 2941 29595 2975
rect 31125 2941 31159 2975
rect 31953 2941 31987 2975
rect 33425 2941 33459 2975
rect 33609 2941 33643 2975
rect 34529 2941 34563 2975
rect 34713 2941 34747 2975
rect 34989 2941 35023 2975
rect 37473 2941 37507 2975
rect 37749 2941 37783 2975
rect 40049 2941 40083 2975
rect 41981 2941 42015 2975
rect 43453 2941 43487 2975
rect 45569 2941 45603 2975
rect 18245 2873 18279 2907
rect 19533 2873 19567 2907
rect 40693 2873 40727 2907
rect 44097 2873 44131 2907
rect 46213 2873 46247 2907
rect 47501 2873 47535 2907
rect 48973 2873 49007 2907
rect 50261 2873 50295 2907
rect 51733 2873 51767 2907
rect 53021 2873 53055 2907
rect 8493 2805 8527 2839
rect 9137 2805 9171 2839
rect 9965 2805 9999 2839
rect 10609 2805 10643 2839
rect 11253 2805 11287 2839
rect 11713 2805 11747 2839
rect 12725 2805 12759 2839
rect 13369 2805 13403 2839
rect 14013 2805 14047 2839
rect 14657 2805 14691 2839
rect 15485 2805 15519 2839
rect 16129 2805 16163 2839
rect 16773 2805 16807 2839
rect 18889 2805 18923 2839
rect 21557 2805 21591 2839
rect 22937 2805 22971 2839
rect 42809 2805 42843 2839
rect 44741 2805 44775 2839
rect 46857 2805 46891 2839
rect 48329 2805 48363 2839
rect 49617 2805 49651 2839
rect 51089 2805 51123 2839
rect 52377 2805 52411 2839
rect 16773 2601 16807 2635
rect 22293 2601 22327 2635
rect 22937 2601 22971 2635
rect 24317 2601 24351 2635
rect 25697 2601 25731 2635
rect 27077 2601 27111 2635
rect 29745 2601 29779 2635
rect 30665 2601 30699 2635
rect 32597 2601 32631 2635
rect 33241 2601 33275 2635
rect 33885 2601 33919 2635
rect 34529 2601 34563 2635
rect 35265 2601 35299 2635
rect 36001 2601 36035 2635
rect 37381 2601 37415 2635
rect 38025 2601 38059 2635
rect 38669 2601 38703 2635
rect 39313 2601 39347 2635
rect 40049 2601 40083 2635
rect 48973 2601 49007 2635
rect 51733 2601 51767 2635
rect 9873 2533 9907 2567
rect 11253 2533 11287 2567
rect 12633 2533 12667 2567
rect 14013 2533 14047 2567
rect 16037 2533 16071 2567
rect 18797 2533 18831 2567
rect 23581 2533 23615 2567
rect 26341 2533 26375 2567
rect 27721 2533 27755 2567
rect 31953 2533 31987 2567
rect 36553 2533 36587 2567
rect 42073 2533 42107 2567
rect 44189 2533 44223 2567
rect 46949 2533 46983 2567
rect 49709 2533 49743 2567
rect 53113 2533 53147 2567
rect 15393 2465 15427 2499
rect 17417 2465 17451 2499
rect 20177 2465 20211 2499
rect 21557 2465 21591 2499
rect 24961 2465 24995 2499
rect 29193 2465 29227 2499
rect 40693 2465 40727 2499
rect 43453 2465 43487 2499
rect 45569 2465 45603 2499
rect 48329 2465 48363 2499
rect 51089 2465 51123 2499
rect 53849 2465 53883 2499
rect 7113 2397 7147 2431
rect 7757 2397 7791 2431
rect 8493 2397 8527 2431
rect 9137 2397 9171 2431
rect 10517 2397 10551 2431
rect 11897 2397 11931 2431
rect 13277 2397 13311 2431
rect 14657 2397 14691 2431
rect 18153 2397 18187 2431
rect 19533 2397 19567 2431
rect 20913 2397 20947 2431
rect 23489 2397 23523 2431
rect 25053 2397 25087 2431
rect 26249 2397 26283 2431
rect 27629 2397 27663 2431
rect 28273 2397 28307 2431
rect 29653 2397 29687 2431
rect 33333 2397 33367 2431
rect 33977 2397 34011 2431
rect 35357 2397 35391 2431
rect 35909 2397 35943 2431
rect 37289 2397 37323 2431
rect 37933 2397 37967 2431
rect 41429 2397 41463 2431
rect 42809 2397 42843 2431
rect 44833 2397 44867 2431
rect 46213 2397 46247 2431
rect 47593 2397 47627 2431
rect 50353 2397 50387 2431
rect 52469 2397 52503 2431
rect 28365 2329 28399 2363
<< metal1 >>
rect 20162 57876 20168 57928
rect 20220 57916 20226 57928
rect 25406 57916 25412 57928
rect 20220 57888 25412 57916
rect 20220 57876 20226 57888
rect 25406 57876 25412 57888
rect 25464 57876 25470 57928
rect 27706 57876 27712 57928
rect 27764 57916 27770 57928
rect 34698 57916 34704 57928
rect 27764 57888 34704 57916
rect 27764 57876 27770 57888
rect 34698 57876 34704 57888
rect 34756 57876 34762 57928
rect 39114 57876 39120 57928
rect 39172 57916 39178 57928
rect 43438 57916 43444 57928
rect 39172 57888 43444 57916
rect 39172 57876 39178 57888
rect 43438 57876 43444 57888
rect 43496 57876 43502 57928
rect 21818 57808 21824 57860
rect 21876 57848 21882 57860
rect 26418 57848 26424 57860
rect 21876 57820 26424 57848
rect 21876 57808 21882 57820
rect 26418 57808 26424 57820
rect 26476 57808 26482 57860
rect 28074 57808 28080 57860
rect 28132 57848 28138 57860
rect 36170 57848 36176 57860
rect 28132 57820 36176 57848
rect 28132 57808 28138 57820
rect 36170 57808 36176 57820
rect 36228 57808 36234 57860
rect 40126 57808 40132 57860
rect 40184 57848 40190 57860
rect 51258 57848 51264 57860
rect 40184 57820 51264 57848
rect 40184 57808 40190 57820
rect 51258 57808 51264 57820
rect 51316 57808 51322 57860
rect 13262 57740 13268 57792
rect 13320 57780 13326 57792
rect 24210 57780 24216 57792
rect 13320 57752 24216 57780
rect 13320 57740 13326 57752
rect 24210 57740 24216 57752
rect 24268 57740 24274 57792
rect 24486 57740 24492 57792
rect 24544 57780 24550 57792
rect 39942 57780 39948 57792
rect 24544 57752 39948 57780
rect 24544 57740 24550 57752
rect 39942 57740 39948 57752
rect 40000 57740 40006 57792
rect 40494 57740 40500 57792
rect 40552 57780 40558 57792
rect 44818 57780 44824 57792
rect 40552 57752 44824 57780
rect 40552 57740 40558 57752
rect 44818 57740 44824 57752
rect 44876 57740 44882 57792
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 3605 57579 3663 57585
rect 3605 57545 3617 57579
rect 3651 57576 3663 57579
rect 3694 57576 3700 57588
rect 3651 57548 3700 57576
rect 3651 57545 3663 57548
rect 3605 57539 3663 57545
rect 3694 57536 3700 57548
rect 3752 57576 3758 57588
rect 3752 57548 4292 57576
rect 3752 57536 3758 57548
rect 4264 57517 4292 57548
rect 5534 57536 5540 57588
rect 5592 57576 5598 57588
rect 5629 57579 5687 57585
rect 5629 57576 5641 57579
rect 5592 57548 5641 57576
rect 5592 57536 5598 57548
rect 5629 57545 5641 57548
rect 5675 57545 5687 57579
rect 5629 57539 5687 57545
rect 10321 57579 10379 57585
rect 10321 57545 10333 57579
rect 10367 57576 10379 57579
rect 10594 57576 10600 57588
rect 10367 57548 10600 57576
rect 10367 57545 10379 57548
rect 10321 57539 10379 57545
rect 10594 57536 10600 57548
rect 10652 57536 10658 57588
rect 11701 57579 11759 57585
rect 11701 57545 11713 57579
rect 11747 57576 11759 57579
rect 11974 57576 11980 57588
rect 11747 57548 11980 57576
rect 11747 57545 11759 57548
rect 11701 57539 11759 57545
rect 11974 57536 11980 57548
rect 12032 57536 12038 57588
rect 13081 57579 13139 57585
rect 13081 57545 13093 57579
rect 13127 57576 13139 57579
rect 13354 57576 13360 57588
rect 13127 57548 13360 57576
rect 13127 57545 13139 57548
rect 13081 57539 13139 57545
rect 13354 57536 13360 57548
rect 13412 57536 13418 57588
rect 14461 57579 14519 57585
rect 14461 57545 14473 57579
rect 14507 57576 14519 57579
rect 14734 57576 14740 57588
rect 14507 57548 14740 57576
rect 14507 57545 14519 57548
rect 14461 57539 14519 57545
rect 14734 57536 14740 57548
rect 14792 57536 14798 57588
rect 15841 57579 15899 57585
rect 15841 57545 15853 57579
rect 15887 57576 15899 57579
rect 16114 57576 16120 57588
rect 15887 57548 16120 57576
rect 15887 57545 15899 57548
rect 15841 57539 15899 57545
rect 16114 57536 16120 57548
rect 16172 57536 16178 57588
rect 17221 57579 17279 57585
rect 17221 57545 17233 57579
rect 17267 57576 17279 57579
rect 17494 57576 17500 57588
rect 17267 57548 17500 57576
rect 17267 57545 17279 57548
rect 17221 57539 17279 57545
rect 17494 57536 17500 57548
rect 17552 57536 17558 57588
rect 18601 57579 18659 57585
rect 18601 57545 18613 57579
rect 18647 57576 18659 57579
rect 18874 57576 18880 57588
rect 18647 57548 18880 57576
rect 18647 57545 18659 57548
rect 18601 57539 18659 57545
rect 18874 57536 18880 57548
rect 18932 57536 18938 57588
rect 19981 57579 20039 57585
rect 19981 57545 19993 57579
rect 20027 57576 20039 57579
rect 20254 57576 20260 57588
rect 20027 57548 20260 57576
rect 20027 57545 20039 57548
rect 19981 57539 20039 57545
rect 20254 57536 20260 57548
rect 20312 57536 20318 57588
rect 21361 57579 21419 57585
rect 21361 57545 21373 57579
rect 21407 57576 21419 57579
rect 21542 57576 21548 57588
rect 21407 57548 21548 57576
rect 21407 57545 21419 57548
rect 21361 57539 21419 57545
rect 21542 57536 21548 57548
rect 21600 57536 21606 57588
rect 22741 57579 22799 57585
rect 22741 57545 22753 57579
rect 22787 57576 22799 57579
rect 24394 57576 24400 57588
rect 22787 57548 24400 57576
rect 22787 57545 22799 57548
rect 22741 57539 22799 57545
rect 24394 57536 24400 57548
rect 24452 57536 24458 57588
rect 28994 57536 29000 57588
rect 29052 57576 29058 57588
rect 29089 57579 29147 57585
rect 29089 57576 29101 57579
rect 29052 57548 29101 57576
rect 29052 57536 29058 57548
rect 29089 57545 29101 57548
rect 29135 57545 29147 57579
rect 29089 57539 29147 57545
rect 29638 57536 29644 57588
rect 29696 57576 29702 57588
rect 29825 57579 29883 57585
rect 29825 57576 29837 57579
rect 29696 57548 29837 57576
rect 29696 57536 29702 57548
rect 29825 57545 29837 57548
rect 29871 57576 29883 57579
rect 30282 57576 30288 57588
rect 29871 57548 30288 57576
rect 29871 57545 29883 57548
rect 29825 57539 29883 57545
rect 30282 57536 30288 57548
rect 30340 57536 30346 57588
rect 30561 57579 30619 57585
rect 30561 57545 30573 57579
rect 30607 57545 30619 57579
rect 30561 57539 30619 57545
rect 4249 57511 4307 57517
rect 4249 57477 4261 57511
rect 4295 57477 4307 57511
rect 21450 57508 21456 57520
rect 4249 57471 4307 57477
rect 16546 57480 21456 57508
rect 5813 57443 5871 57449
rect 5813 57409 5825 57443
rect 5859 57440 5871 57443
rect 6362 57440 6368 57452
rect 5859 57412 6368 57440
rect 5859 57409 5871 57412
rect 5813 57403 5871 57409
rect 6362 57400 6368 57412
rect 6420 57400 6426 57452
rect 7374 57400 7380 57452
rect 7432 57440 7438 57452
rect 7469 57443 7527 57449
rect 7469 57440 7481 57443
rect 7432 57412 7481 57440
rect 7432 57400 7438 57412
rect 7469 57409 7481 57412
rect 7515 57409 7527 57443
rect 8294 57440 8300 57452
rect 8255 57412 8300 57440
rect 7469 57403 7527 57409
rect 8294 57400 8300 57412
rect 8352 57400 8358 57452
rect 9125 57443 9183 57449
rect 9125 57409 9137 57443
rect 9171 57440 9183 57443
rect 9214 57440 9220 57452
rect 9171 57412 9220 57440
rect 9171 57409 9183 57412
rect 9125 57403 9183 57409
rect 9214 57400 9220 57412
rect 9272 57400 9278 57452
rect 10505 57443 10563 57449
rect 10505 57409 10517 57443
rect 10551 57440 10563 57443
rect 11882 57440 11888 57452
rect 10551 57412 11192 57440
rect 11843 57412 11888 57440
rect 10551 57409 10563 57412
rect 10505 57403 10563 57409
rect 4433 57307 4491 57313
rect 4433 57273 4445 57307
rect 4479 57304 4491 57307
rect 11054 57304 11060 57316
rect 4479 57276 11060 57304
rect 4479 57273 4491 57276
rect 4433 57267 4491 57273
rect 11054 57264 11060 57276
rect 11112 57264 11118 57316
rect 11164 57245 11192 57412
rect 11882 57400 11888 57412
rect 11940 57400 11946 57452
rect 13262 57440 13268 57452
rect 13223 57412 13268 57440
rect 13262 57400 13268 57412
rect 13320 57400 13326 57452
rect 14645 57443 14703 57449
rect 14645 57409 14657 57443
rect 14691 57409 14703 57443
rect 14645 57403 14703 57409
rect 16025 57443 16083 57449
rect 16025 57409 16037 57443
rect 16071 57440 16083 57443
rect 16546 57440 16574 57480
rect 21450 57468 21456 57480
rect 21508 57468 21514 57520
rect 21726 57468 21732 57520
rect 21784 57508 21790 57520
rect 26970 57508 26976 57520
rect 21784 57480 26976 57508
rect 21784 57468 21790 57480
rect 26970 57468 26976 57480
rect 27028 57468 27034 57520
rect 27154 57468 27160 57520
rect 27212 57508 27218 57520
rect 27212 57480 28028 57508
rect 27212 57468 27218 57480
rect 17402 57440 17408 57452
rect 16071 57412 16574 57440
rect 17363 57412 17408 57440
rect 16071 57409 16083 57412
rect 16025 57403 16083 57409
rect 14660 57304 14688 57403
rect 17402 57400 17408 57412
rect 17460 57400 17466 57452
rect 18785 57443 18843 57449
rect 18785 57409 18797 57443
rect 18831 57409 18843 57443
rect 20162 57440 20168 57452
rect 20123 57412 20168 57440
rect 18785 57403 18843 57409
rect 18800 57372 18828 57403
rect 20162 57400 20168 57412
rect 20220 57400 20226 57452
rect 21545 57443 21603 57449
rect 21545 57409 21557 57443
rect 21591 57438 21603 57443
rect 21818 57440 21824 57452
rect 21652 57438 21824 57440
rect 21591 57412 21824 57438
rect 21591 57410 21680 57412
rect 21591 57409 21603 57410
rect 21545 57403 21603 57409
rect 21818 57400 21824 57412
rect 21876 57400 21882 57452
rect 21910 57400 21916 57452
rect 21968 57440 21974 57452
rect 22925 57443 22983 57449
rect 21968 57412 22876 57440
rect 21968 57400 21974 57412
rect 22278 57372 22284 57384
rect 18800 57344 22284 57372
rect 22278 57332 22284 57344
rect 22336 57332 22342 57384
rect 22848 57372 22876 57412
rect 22925 57409 22937 57443
rect 22971 57440 22983 57443
rect 23750 57440 23756 57452
rect 22971 57412 23756 57440
rect 22971 57409 22983 57412
rect 22925 57403 22983 57409
rect 23750 57400 23756 57412
rect 23808 57400 23814 57452
rect 24118 57440 24124 57452
rect 24079 57412 24124 57440
rect 24118 57400 24124 57412
rect 24176 57400 24182 57452
rect 24302 57440 24308 57452
rect 24263 57412 24308 57440
rect 24302 57400 24308 57412
rect 24360 57400 24366 57452
rect 25222 57400 25228 57452
rect 25280 57440 25286 57452
rect 25317 57443 25375 57449
rect 25317 57440 25329 57443
rect 25280 57412 25329 57440
rect 25280 57400 25286 57412
rect 25317 57409 25329 57412
rect 25363 57409 25375 57443
rect 25498 57440 25504 57452
rect 25411 57412 25504 57440
rect 25317 57403 25375 57409
rect 25498 57400 25504 57412
rect 25556 57440 25562 57452
rect 25556 57412 26832 57440
rect 25556 57400 25562 57412
rect 23658 57372 23664 57384
rect 22848 57344 23664 57372
rect 23658 57332 23664 57344
rect 23716 57372 23722 57384
rect 23937 57375 23995 57381
rect 23937 57372 23949 57375
rect 23716 57344 23949 57372
rect 23716 57332 23722 57344
rect 23937 57341 23949 57344
rect 23983 57341 23995 57375
rect 26234 57372 26240 57384
rect 23937 57335 23995 57341
rect 25516 57344 26240 57372
rect 25038 57304 25044 57316
rect 14660 57276 25044 57304
rect 25038 57264 25044 57276
rect 25096 57264 25102 57316
rect 11149 57239 11207 57245
rect 11149 57205 11161 57239
rect 11195 57236 11207 57239
rect 20714 57236 20720 57248
rect 11195 57208 20720 57236
rect 11195 57205 11207 57208
rect 11149 57199 11207 57205
rect 20714 57196 20720 57208
rect 20772 57196 20778 57248
rect 20809 57239 20867 57245
rect 20809 57205 20821 57239
rect 20855 57236 20867 57239
rect 21910 57236 21916 57248
rect 20855 57208 21916 57236
rect 20855 57205 20867 57208
rect 20809 57199 20867 57205
rect 21910 57196 21916 57208
rect 21968 57196 21974 57248
rect 22094 57236 22100 57248
rect 22055 57208 22100 57236
rect 22094 57196 22100 57208
rect 22152 57236 22158 57248
rect 25516 57236 25544 57344
rect 26234 57332 26240 57344
rect 26292 57372 26298 57384
rect 26697 57375 26755 57381
rect 26697 57372 26709 57375
rect 26292 57344 26709 57372
rect 26292 57332 26298 57344
rect 26697 57341 26709 57344
rect 26743 57341 26755 57375
rect 26697 57335 26755 57341
rect 26804 57304 26832 57412
rect 26878 57400 26884 57452
rect 26936 57440 26942 57452
rect 27706 57440 27712 57452
rect 26936 57412 26981 57440
rect 27632 57412 27712 57440
rect 26936 57400 26942 57412
rect 27632 57384 27660 57412
rect 27706 57400 27712 57412
rect 27764 57400 27770 57452
rect 27890 57440 27896 57452
rect 27851 57412 27896 57440
rect 27890 57400 27896 57412
rect 27948 57400 27954 57452
rect 28000 57440 28028 57480
rect 28166 57468 28172 57520
rect 28224 57508 28230 57520
rect 30576 57508 30604 57539
rect 30650 57536 30656 57588
rect 30708 57576 30714 57588
rect 35526 57576 35532 57588
rect 30708 57548 35532 57576
rect 30708 57536 30714 57548
rect 35526 57536 35532 57548
rect 35584 57536 35590 57588
rect 39942 57536 39948 57588
rect 40000 57576 40006 57588
rect 40037 57579 40095 57585
rect 40037 57576 40049 57579
rect 40000 57548 40049 57576
rect 40000 57536 40006 57548
rect 40037 57545 40049 57548
rect 40083 57545 40095 57579
rect 40037 57539 40095 57545
rect 42153 57579 42211 57585
rect 42153 57545 42165 57579
rect 42199 57576 42211 57579
rect 43806 57576 43812 57588
rect 42199 57548 43812 57576
rect 42199 57545 42211 57548
rect 42153 57539 42211 57545
rect 43806 57536 43812 57548
rect 43864 57536 43870 57588
rect 43990 57536 43996 57588
rect 44048 57576 44054 57588
rect 51258 57576 51264 57588
rect 44048 57548 48636 57576
rect 51219 57548 51264 57576
rect 44048 57536 44054 57548
rect 28224 57480 30604 57508
rect 28224 57468 28230 57480
rect 32950 57468 32956 57520
rect 33008 57508 33014 57520
rect 33008 57480 34744 57508
rect 33008 57468 33014 57480
rect 29273 57443 29331 57449
rect 28000 57412 28994 57440
rect 27614 57372 27620 57384
rect 27527 57344 27620 57372
rect 27614 57332 27620 57344
rect 27672 57332 27678 57384
rect 28166 57372 28172 57384
rect 27724 57344 28172 57372
rect 27724 57304 27752 57344
rect 28166 57332 28172 57344
rect 28224 57332 28230 57384
rect 28966 57372 28994 57412
rect 29273 57409 29285 57443
rect 29319 57440 29331 57443
rect 29454 57440 29460 57452
rect 29319 57412 29460 57440
rect 29319 57409 29331 57412
rect 29273 57403 29331 57409
rect 29454 57400 29460 57412
rect 29512 57400 29518 57452
rect 30377 57443 30435 57449
rect 30377 57409 30389 57443
rect 30423 57409 30435 57443
rect 30377 57403 30435 57409
rect 30392 57372 30420 57403
rect 31754 57400 31760 57452
rect 31812 57440 31818 57452
rect 33321 57443 33379 57449
rect 31812 57412 31857 57440
rect 31812 57400 31818 57412
rect 33321 57409 33333 57443
rect 33367 57440 33379 57443
rect 33686 57440 33692 57452
rect 33367 57412 33692 57440
rect 33367 57409 33379 57412
rect 33321 57403 33379 57409
rect 33686 57400 33692 57412
rect 33744 57400 33750 57452
rect 33778 57400 33784 57452
rect 33836 57440 33842 57452
rect 34716 57449 34744 57480
rect 35618 57468 35624 57520
rect 35676 57508 35682 57520
rect 35676 57480 37596 57508
rect 35676 57468 35682 57480
rect 34517 57443 34575 57449
rect 34517 57440 34529 57443
rect 33836 57412 34529 57440
rect 33836 57400 33842 57412
rect 34517 57409 34529 57412
rect 34563 57409 34575 57443
rect 34517 57403 34575 57409
rect 34701 57443 34759 57449
rect 34701 57409 34713 57443
rect 34747 57409 34759 57443
rect 34701 57403 34759 57409
rect 34790 57400 34796 57452
rect 34848 57440 34854 57452
rect 34977 57443 35035 57449
rect 34977 57440 34989 57443
rect 34848 57412 34989 57440
rect 34848 57400 34854 57412
rect 34977 57409 34989 57412
rect 35023 57440 35035 57443
rect 36173 57443 36231 57449
rect 36173 57440 36185 57443
rect 35023 57412 36185 57440
rect 35023 57409 35035 57412
rect 34977 57403 35035 57409
rect 36173 57409 36185 57412
rect 36219 57440 36231 57443
rect 36262 57440 36268 57452
rect 36219 57412 36268 57440
rect 36219 57409 36231 57412
rect 36173 57403 36231 57409
rect 36262 57400 36268 57412
rect 36320 57400 36326 57452
rect 37568 57449 37596 57480
rect 40218 57468 40224 57520
rect 40276 57508 40282 57520
rect 44008 57508 44036 57536
rect 40276 57480 40448 57508
rect 40276 57468 40282 57480
rect 37553 57443 37611 57449
rect 37553 57409 37565 57443
rect 37599 57409 37611 57443
rect 38654 57440 38660 57452
rect 38567 57412 38660 57440
rect 37553 57403 37611 57409
rect 38654 57400 38660 57412
rect 38712 57440 38718 57452
rect 39850 57440 39856 57452
rect 38712 57412 39856 57440
rect 38712 57400 38718 57412
rect 39850 57400 39856 57412
rect 39908 57400 39914 57452
rect 40420 57449 40448 57480
rect 41984 57480 44036 57508
rect 41984 57449 42012 57480
rect 45554 57468 45560 57520
rect 45612 57508 45618 57520
rect 45830 57508 45836 57520
rect 45612 57480 45836 57508
rect 45612 57468 45618 57480
rect 45830 57468 45836 57480
rect 45888 57468 45894 57520
rect 40405 57443 40463 57449
rect 40405 57409 40417 57443
rect 40451 57409 40463 57443
rect 40405 57403 40463 57409
rect 41969 57443 42027 57449
rect 41969 57409 41981 57443
rect 42015 57409 42027 57443
rect 41969 57403 42027 57409
rect 42245 57443 42303 57449
rect 42245 57409 42257 57443
rect 42291 57440 42303 57443
rect 44361 57443 44419 57449
rect 42291 57412 43116 57440
rect 42291 57409 42303 57412
rect 42245 57403 42303 57409
rect 43088 57384 43116 57412
rect 44361 57409 44373 57443
rect 44407 57409 44419 57443
rect 46934 57440 46940 57452
rect 46895 57412 46940 57440
rect 44361 57403 44419 57409
rect 28966 57344 30420 57372
rect 32033 57375 32091 57381
rect 32033 57341 32045 57375
rect 32079 57372 32091 57375
rect 32398 57372 32404 57384
rect 32079 57344 32404 57372
rect 32079 57341 32091 57344
rect 32033 57335 32091 57341
rect 32398 57332 32404 57344
rect 32456 57332 32462 57384
rect 33597 57375 33655 57381
rect 33597 57341 33609 57375
rect 33643 57372 33655 57375
rect 35894 57372 35900 57384
rect 33643 57344 34652 57372
rect 35855 57344 35900 57372
rect 33643 57341 33655 57344
rect 33597 57335 33655 57341
rect 34624 57316 34652 57344
rect 35894 57332 35900 57344
rect 35952 57332 35958 57384
rect 37274 57372 37280 57384
rect 37187 57344 37280 57372
rect 37274 57332 37280 57344
rect 37332 57372 37338 57384
rect 37458 57372 37464 57384
rect 37332 57344 37464 57372
rect 37332 57332 37338 57344
rect 37458 57332 37464 57344
rect 37516 57332 37522 57384
rect 38933 57375 38991 57381
rect 38933 57341 38945 57375
rect 38979 57341 38991 57375
rect 38933 57335 38991 57341
rect 40221 57375 40279 57381
rect 40221 57341 40233 57375
rect 40267 57341 40279 57375
rect 40221 57335 40279 57341
rect 26804 57276 27752 57304
rect 27801 57307 27859 57313
rect 27801 57273 27813 57307
rect 27847 57304 27859 57307
rect 28258 57304 28264 57316
rect 27847 57276 28264 57304
rect 27847 57273 27859 57276
rect 27801 57267 27859 57273
rect 28258 57264 28264 57276
rect 28316 57264 28322 57316
rect 28902 57264 28908 57316
rect 28960 57304 28966 57316
rect 33137 57307 33195 57313
rect 33137 57304 33149 57307
rect 28960 57276 33149 57304
rect 28960 57264 28966 57276
rect 33137 57273 33149 57276
rect 33183 57273 33195 57307
rect 33137 57267 33195 57273
rect 33410 57264 33416 57316
rect 33468 57304 33474 57316
rect 33505 57307 33563 57313
rect 33505 57304 33517 57307
rect 33468 57276 33517 57304
rect 33468 57264 33474 57276
rect 33505 57273 33517 57276
rect 33551 57304 33563 57307
rect 33551 57276 34560 57304
rect 33551 57273 33563 57276
rect 33505 57267 33563 57273
rect 22152 57208 25544 57236
rect 22152 57196 22158 57208
rect 25590 57196 25596 57248
rect 25648 57236 25654 57248
rect 25685 57239 25743 57245
rect 25685 57236 25697 57239
rect 25648 57208 25697 57236
rect 25648 57196 25654 57208
rect 25685 57205 25697 57208
rect 25731 57205 25743 57239
rect 27062 57236 27068 57248
rect 27023 57208 27068 57236
rect 25685 57199 25743 57205
rect 27062 57196 27068 57208
rect 27120 57196 27126 57248
rect 27706 57236 27712 57248
rect 27667 57208 27712 57236
rect 27706 57196 27712 57208
rect 27764 57196 27770 57248
rect 28445 57239 28503 57245
rect 28445 57205 28457 57239
rect 28491 57236 28503 57239
rect 29270 57236 29276 57248
rect 28491 57208 29276 57236
rect 28491 57205 28503 57208
rect 28445 57199 28503 57205
rect 29270 57196 29276 57208
rect 29328 57196 29334 57248
rect 29362 57196 29368 57248
rect 29420 57236 29426 57248
rect 30650 57236 30656 57248
rect 29420 57208 30656 57236
rect 29420 57196 29426 57208
rect 30650 57196 30656 57208
rect 30708 57196 30714 57248
rect 31018 57196 31024 57248
rect 31076 57236 31082 57248
rect 31113 57239 31171 57245
rect 31113 57236 31125 57239
rect 31076 57208 31125 57236
rect 31076 57196 31082 57208
rect 31113 57205 31125 57208
rect 31159 57205 31171 57239
rect 31113 57199 31171 57205
rect 32214 57196 32220 57248
rect 32272 57236 32278 57248
rect 34330 57236 34336 57248
rect 32272 57208 34336 57236
rect 32272 57196 32278 57208
rect 34330 57196 34336 57208
rect 34388 57196 34394 57248
rect 34532 57236 34560 57276
rect 34606 57264 34612 57316
rect 34664 57304 34670 57316
rect 38948 57304 38976 57335
rect 34664 57276 38976 57304
rect 40236 57304 40264 57335
rect 40310 57332 40316 57384
rect 40368 57372 40374 57384
rect 40368 57344 40413 57372
rect 40368 57332 40374 57344
rect 40494 57332 40500 57384
rect 40552 57372 40558 57384
rect 42797 57375 42855 57381
rect 40552 57344 40597 57372
rect 40552 57332 40558 57344
rect 42797 57341 42809 57375
rect 42843 57372 42855 57375
rect 42886 57372 42892 57384
rect 42843 57344 42892 57372
rect 42843 57341 42855 57344
rect 42797 57335 42855 57341
rect 42886 57332 42892 57344
rect 42944 57332 42950 57384
rect 43070 57372 43076 57384
rect 43031 57344 43076 57372
rect 43070 57332 43076 57344
rect 43128 57332 43134 57384
rect 43806 57332 43812 57384
rect 43864 57372 43870 57384
rect 44376 57372 44404 57403
rect 46934 57400 46940 57412
rect 46992 57400 46998 57452
rect 48314 57440 48320 57452
rect 48275 57412 48320 57440
rect 48314 57400 48320 57412
rect 48372 57400 48378 57452
rect 48608 57449 48636 57548
rect 51258 57536 51264 57548
rect 51316 57536 51322 57588
rect 52454 57536 52460 57588
rect 52512 57536 52518 57588
rect 52472 57508 52500 57536
rect 52546 57508 52552 57520
rect 52459 57480 52552 57508
rect 52546 57468 52552 57480
rect 52604 57508 52610 57520
rect 52641 57511 52699 57517
rect 52641 57508 52653 57511
rect 52604 57480 52653 57508
rect 52604 57468 52610 57480
rect 52641 57477 52653 57480
rect 52687 57477 52699 57511
rect 52641 57471 52699 57477
rect 48593 57443 48651 57449
rect 48593 57409 48605 57443
rect 48639 57409 48651 57443
rect 49694 57440 49700 57452
rect 49655 57412 49700 57440
rect 48593 57403 48651 57409
rect 49694 57400 49700 57412
rect 49752 57400 49758 57452
rect 51074 57400 51080 57452
rect 51132 57440 51138 57452
rect 51445 57443 51503 57449
rect 51445 57440 51457 57443
rect 51132 57412 51457 57440
rect 51132 57400 51138 57412
rect 51445 57409 51457 57412
rect 51491 57440 51503 57443
rect 51626 57440 51632 57452
rect 51491 57412 51632 57440
rect 51491 57409 51503 57412
rect 51445 57403 51503 57409
rect 51626 57400 51632 57412
rect 51684 57400 51690 57452
rect 53834 57400 53840 57452
rect 53892 57440 53898 57452
rect 53929 57443 53987 57449
rect 53929 57440 53941 57443
rect 53892 57412 53941 57440
rect 53892 57400 53898 57412
rect 53929 57409 53941 57412
rect 53975 57409 53987 57443
rect 53929 57403 53987 57409
rect 55214 57400 55220 57452
rect 55272 57440 55278 57452
rect 55309 57443 55367 57449
rect 55309 57440 55321 57443
rect 55272 57412 55321 57440
rect 55272 57400 55278 57412
rect 55309 57409 55321 57412
rect 55355 57409 55367 57443
rect 55309 57403 55367 57409
rect 55674 57400 55680 57452
rect 55732 57440 55738 57452
rect 56597 57443 56655 57449
rect 56597 57440 56609 57443
rect 55732 57412 56609 57440
rect 55732 57400 55738 57412
rect 56597 57409 56609 57412
rect 56643 57409 56655 57443
rect 56597 57403 56655 57409
rect 44542 57372 44548 57384
rect 43864 57344 44312 57372
rect 44376 57344 44548 57372
rect 43864 57332 43870 57344
rect 40586 57304 40592 57316
rect 40236 57276 40592 57304
rect 34664 57264 34670 57276
rect 40586 57264 40592 57276
rect 40644 57264 40650 57316
rect 34885 57239 34943 57245
rect 34885 57236 34897 57239
rect 34532 57208 34897 57236
rect 34885 57205 34897 57208
rect 34931 57236 34943 57239
rect 36446 57236 36452 57248
rect 34931 57208 36452 57236
rect 34931 57205 34943 57208
rect 34885 57199 34943 57205
rect 36446 57196 36452 57208
rect 36504 57236 36510 57248
rect 40126 57236 40132 57248
rect 36504 57208 40132 57236
rect 36504 57196 36510 57208
rect 40126 57196 40132 57208
rect 40184 57196 40190 57248
rect 40770 57196 40776 57248
rect 40828 57236 40834 57248
rect 41785 57239 41843 57245
rect 41785 57236 41797 57239
rect 40828 57208 41797 57236
rect 40828 57196 40834 57208
rect 41785 57205 41797 57208
rect 41831 57205 41843 57239
rect 44174 57236 44180 57248
rect 44135 57208 44180 57236
rect 41785 57199 41843 57205
rect 44174 57196 44180 57208
rect 44232 57196 44238 57248
rect 44284 57236 44312 57344
rect 44542 57332 44548 57344
rect 44600 57332 44606 57384
rect 44637 57375 44695 57381
rect 44637 57341 44649 57375
rect 44683 57372 44695 57375
rect 44726 57372 44732 57384
rect 44683 57344 44732 57372
rect 44683 57341 44695 57344
rect 44637 57335 44695 57341
rect 44726 57332 44732 57344
rect 44784 57372 44790 57384
rect 47210 57372 47216 57384
rect 44784 57344 45600 57372
rect 47171 57344 47216 57372
rect 44784 57332 44790 57344
rect 45572 57304 45600 57344
rect 47210 57332 47216 57344
rect 47268 57332 47274 57384
rect 49973 57375 50031 57381
rect 49973 57341 49985 57375
rect 50019 57341 50031 57375
rect 49973 57335 50031 57341
rect 49988 57304 50016 57335
rect 45572 57276 50016 57304
rect 50062 57264 50068 57316
rect 50120 57304 50126 57316
rect 55493 57307 55551 57313
rect 55493 57304 55505 57307
rect 50120 57276 55505 57304
rect 50120 57264 50126 57276
rect 55493 57273 55505 57276
rect 55539 57273 55551 57307
rect 55493 57267 55551 57273
rect 44545 57239 44603 57245
rect 44545 57236 44557 57239
rect 44284 57208 44557 57236
rect 44545 57205 44557 57208
rect 44591 57236 44603 57239
rect 45002 57236 45008 57248
rect 44591 57208 45008 57236
rect 44591 57205 44603 57208
rect 44545 57199 44603 57205
rect 45002 57196 45008 57208
rect 45060 57196 45066 57248
rect 45738 57236 45744 57248
rect 45699 57208 45744 57236
rect 45738 57196 45744 57208
rect 45796 57196 45802 57248
rect 51074 57196 51080 57248
rect 51132 57236 51138 57248
rect 52733 57239 52791 57245
rect 52733 57236 52745 57239
rect 51132 57208 52745 57236
rect 51132 57196 51138 57208
rect 52733 57205 52745 57208
rect 52779 57205 52791 57239
rect 54110 57236 54116 57248
rect 54071 57208 54116 57236
rect 52733 57199 52791 57205
rect 54110 57196 54116 57208
rect 54168 57196 54174 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 4614 56992 4620 57044
rect 4672 57032 4678 57044
rect 4709 57035 4767 57041
rect 4709 57032 4721 57035
rect 4672 57004 4721 57032
rect 4672 56992 4678 57004
rect 4709 57001 4721 57004
rect 4755 57001 4767 57035
rect 4709 56995 4767 57001
rect 5905 57035 5963 57041
rect 5905 57001 5917 57035
rect 5951 57032 5963 57035
rect 5994 57032 6000 57044
rect 5951 57004 6000 57032
rect 5951 57001 5963 57004
rect 5905 56995 5963 57001
rect 5994 56992 6000 57004
rect 6052 56992 6058 57044
rect 6454 56992 6460 57044
rect 6512 57032 6518 57044
rect 6549 57035 6607 57041
rect 6549 57032 6561 57035
rect 6512 57004 6561 57032
rect 6512 56992 6518 57004
rect 6549 57001 6561 57004
rect 6595 57001 6607 57035
rect 6549 56995 6607 57001
rect 8754 56992 8760 57044
rect 8812 57032 8818 57044
rect 8849 57035 8907 57041
rect 8849 57032 8861 57035
rect 8812 57004 8861 57032
rect 8812 56992 8818 57004
rect 8849 57001 8861 57004
rect 8895 57001 8907 57035
rect 8849 56995 8907 57001
rect 10134 56992 10140 57044
rect 10192 57032 10198 57044
rect 10229 57035 10287 57041
rect 10229 57032 10241 57035
rect 10192 57004 10241 57032
rect 10192 56992 10198 57004
rect 10229 57001 10241 57004
rect 10275 57001 10287 57035
rect 10229 56995 10287 57001
rect 11514 56992 11520 57044
rect 11572 57032 11578 57044
rect 11609 57035 11667 57041
rect 11609 57032 11621 57035
rect 11572 57004 11621 57032
rect 11572 56992 11578 57004
rect 11609 57001 11621 57004
rect 11655 57001 11667 57035
rect 11609 56995 11667 57001
rect 12894 56992 12900 57044
rect 12952 57032 12958 57044
rect 12989 57035 13047 57041
rect 12989 57032 13001 57035
rect 12952 57004 13001 57032
rect 12952 56992 12958 57004
rect 12989 57001 13001 57004
rect 13035 57001 13047 57035
rect 12989 56995 13047 57001
rect 14274 56992 14280 57044
rect 14332 57032 14338 57044
rect 14369 57035 14427 57041
rect 14369 57032 14381 57035
rect 14332 57004 14381 57032
rect 14332 56992 14338 57004
rect 14369 57001 14381 57004
rect 14415 57001 14427 57035
rect 14369 56995 14427 57001
rect 15654 56992 15660 57044
rect 15712 57032 15718 57044
rect 15749 57035 15807 57041
rect 15749 57032 15761 57035
rect 15712 57004 15761 57032
rect 15712 56992 15718 57004
rect 15749 57001 15761 57004
rect 15795 57001 15807 57035
rect 15749 56995 15807 57001
rect 17034 56992 17040 57044
rect 17092 57032 17098 57044
rect 17129 57035 17187 57041
rect 17129 57032 17141 57035
rect 17092 57004 17141 57032
rect 17092 56992 17098 57004
rect 17129 57001 17141 57004
rect 17175 57001 17187 57035
rect 17129 56995 17187 57001
rect 18414 56992 18420 57044
rect 18472 57032 18478 57044
rect 18509 57035 18567 57041
rect 18509 57032 18521 57035
rect 18472 57004 18521 57032
rect 18472 56992 18478 57004
rect 18509 57001 18521 57004
rect 18555 57001 18567 57035
rect 18509 56995 18567 57001
rect 19889 57035 19947 57041
rect 19889 57001 19901 57035
rect 19935 57032 19947 57035
rect 19978 57032 19984 57044
rect 19935 57004 19984 57032
rect 19935 57001 19947 57004
rect 19889 56995 19947 57001
rect 19978 56992 19984 57004
rect 20036 56992 20042 57044
rect 21174 56992 21180 57044
rect 21232 57032 21238 57044
rect 21269 57035 21327 57041
rect 21269 57032 21281 57035
rect 21232 57004 21281 57032
rect 21232 56992 21238 57004
rect 21269 57001 21281 57004
rect 21315 57001 21327 57035
rect 23014 57032 23020 57044
rect 22975 57004 23020 57032
rect 21269 56995 21327 57001
rect 23014 56992 23020 57004
rect 23072 56992 23078 57044
rect 24210 56992 24216 57044
rect 24268 57032 24274 57044
rect 24305 57035 24363 57041
rect 24305 57032 24317 57035
rect 24268 57004 24317 57032
rect 24268 56992 24274 57004
rect 24305 57001 24317 57004
rect 24351 57001 24363 57035
rect 24305 56995 24363 57001
rect 26970 56992 26976 57044
rect 27028 57032 27034 57044
rect 27065 57035 27123 57041
rect 27065 57032 27077 57035
rect 27028 57004 27077 57032
rect 27028 56992 27034 57004
rect 27065 57001 27077 57004
rect 27111 57001 27123 57035
rect 28074 57032 28080 57044
rect 28035 57004 28080 57032
rect 27065 56995 27123 57001
rect 28074 56992 28080 57004
rect 28132 56992 28138 57044
rect 28166 56992 28172 57044
rect 28224 57032 28230 57044
rect 32674 57032 32680 57044
rect 28224 57004 32680 57032
rect 28224 56992 28230 57004
rect 32674 56992 32680 57004
rect 32732 56992 32738 57044
rect 34241 57035 34299 57041
rect 34241 57032 34253 57035
rect 32784 57004 34253 57032
rect 22278 56964 22284 56976
rect 22191 56936 22284 56964
rect 22278 56924 22284 56936
rect 22336 56924 22342 56976
rect 27617 56967 27675 56973
rect 27617 56933 27629 56967
rect 27663 56964 27675 56967
rect 27982 56964 27988 56976
rect 27663 56936 27988 56964
rect 27663 56933 27675 56936
rect 27617 56927 27675 56933
rect 27982 56924 27988 56936
rect 28040 56924 28046 56976
rect 28442 56924 28448 56976
rect 28500 56964 28506 56976
rect 28902 56964 28908 56976
rect 28500 56936 28908 56964
rect 28500 56924 28506 56936
rect 28902 56924 28908 56936
rect 28960 56964 28966 56976
rect 28960 56936 29316 56964
rect 28960 56924 28966 56936
rect 11054 56856 11060 56908
rect 11112 56896 11118 56908
rect 22094 56896 22100 56908
rect 11112 56868 22100 56896
rect 11112 56856 11118 56868
rect 22094 56856 22100 56868
rect 22152 56856 22158 56908
rect 22296 56896 22324 56924
rect 23661 56899 23719 56905
rect 23661 56896 23673 56899
rect 22296 56868 23673 56896
rect 23661 56865 23673 56868
rect 23707 56865 23719 56899
rect 23661 56859 23719 56865
rect 25406 56856 25412 56908
rect 25464 56896 25470 56908
rect 25685 56899 25743 56905
rect 25464 56868 25636 56896
rect 25464 56856 25470 56868
rect 22465 56831 22523 56837
rect 22465 56797 22477 56831
rect 22511 56797 22523 56831
rect 23198 56828 23204 56840
rect 23159 56800 23204 56828
rect 22465 56791 22523 56797
rect 22480 56760 22508 56791
rect 23198 56788 23204 56800
rect 23256 56788 23262 56840
rect 23750 56828 23756 56840
rect 23711 56800 23756 56828
rect 23750 56788 23756 56800
rect 23808 56788 23814 56840
rect 24118 56828 24124 56840
rect 24090 56800 24124 56828
rect 24118 56788 24124 56800
rect 24176 56837 24182 56840
rect 24176 56831 24238 56837
rect 24176 56797 24192 56831
rect 24226 56828 24238 56831
rect 25314 56831 25372 56837
rect 24226 56800 25268 56828
rect 24226 56797 24238 56800
rect 24176 56791 24238 56797
rect 24176 56788 24182 56791
rect 24026 56760 24032 56772
rect 22480 56732 24032 56760
rect 24026 56720 24032 56732
rect 24084 56720 24090 56772
rect 25240 56760 25268 56800
rect 25314 56797 25326 56831
rect 25360 56828 25372 56831
rect 25498 56828 25504 56840
rect 25360 56800 25504 56828
rect 25360 56797 25372 56800
rect 25314 56791 25372 56797
rect 25498 56788 25504 56800
rect 25556 56788 25562 56840
rect 25608 56828 25636 56868
rect 25685 56865 25697 56899
rect 25731 56896 25743 56899
rect 25866 56896 25872 56908
rect 25731 56868 25872 56896
rect 25731 56865 25743 56868
rect 25685 56859 25743 56865
rect 25866 56856 25872 56868
rect 25924 56856 25930 56908
rect 26418 56896 26424 56908
rect 26379 56868 26424 56896
rect 26418 56856 26424 56868
rect 26476 56856 26482 56908
rect 26510 56856 26516 56908
rect 26568 56896 26574 56908
rect 27154 56896 27160 56908
rect 26568 56868 27160 56896
rect 26568 56856 26574 56868
rect 27154 56856 27160 56868
rect 27212 56856 27218 56908
rect 27706 56856 27712 56908
rect 27764 56896 27770 56908
rect 29178 56896 29184 56908
rect 27764 56868 27936 56896
rect 27764 56856 27770 56868
rect 25777 56831 25835 56837
rect 25777 56828 25789 56831
rect 25608 56800 25789 56828
rect 25777 56797 25789 56800
rect 25823 56797 25835 56831
rect 25777 56791 25835 56797
rect 26940 56831 26998 56837
rect 26940 56797 26952 56831
rect 26986 56828 26998 56831
rect 27338 56828 27344 56840
rect 26986 56800 27344 56828
rect 26986 56797 26998 56800
rect 26940 56791 26998 56797
rect 27338 56788 27344 56800
rect 27396 56788 27402 56840
rect 27430 56788 27436 56840
rect 27488 56828 27494 56840
rect 27908 56837 27936 56868
rect 28000 56868 29184 56896
rect 27801 56831 27859 56837
rect 27801 56828 27813 56831
rect 27488 56800 27813 56828
rect 27488 56788 27494 56800
rect 27801 56797 27813 56800
rect 27847 56797 27859 56831
rect 27801 56791 27859 56797
rect 27893 56831 27951 56837
rect 27893 56797 27905 56831
rect 27939 56797 27951 56831
rect 27893 56791 27951 56797
rect 27522 56760 27528 56772
rect 25240 56732 27528 56760
rect 27522 56720 27528 56732
rect 27580 56720 27586 56772
rect 27816 56760 27844 56791
rect 28000 56760 28028 56868
rect 29178 56856 29184 56868
rect 29236 56856 29242 56908
rect 29288 56896 29316 56936
rect 29362 56924 29368 56976
rect 29420 56964 29426 56976
rect 29546 56964 29552 56976
rect 29420 56936 29552 56964
rect 29420 56924 29426 56936
rect 29546 56924 29552 56936
rect 29604 56924 29610 56976
rect 32784 56964 32812 57004
rect 34241 57001 34253 57004
rect 34287 57001 34299 57035
rect 34241 56995 34299 57001
rect 37277 57035 37335 57041
rect 37277 57001 37289 57035
rect 37323 57032 37335 57035
rect 37366 57032 37372 57044
rect 37323 57004 37372 57032
rect 37323 57001 37335 57004
rect 37277 56995 37335 57001
rect 37366 56992 37372 57004
rect 37424 56992 37430 57044
rect 37568 57004 44312 57032
rect 34790 56964 34796 56976
rect 30944 56936 32812 56964
rect 33704 56936 34796 56964
rect 30944 56896 30972 56936
rect 29288 56868 29684 56896
rect 28166 56828 28172 56840
rect 28127 56800 28172 56828
rect 28166 56788 28172 56800
rect 28224 56788 28230 56840
rect 29270 56828 29276 56840
rect 29231 56800 29276 56828
rect 29270 56788 29276 56800
rect 29328 56788 29334 56840
rect 29362 56788 29368 56840
rect 29420 56828 29426 56840
rect 29656 56837 29684 56868
rect 29932 56868 30972 56896
rect 31113 56899 31171 56905
rect 29457 56831 29515 56837
rect 29457 56828 29469 56831
rect 29420 56800 29469 56828
rect 29420 56788 29426 56800
rect 29457 56797 29469 56800
rect 29503 56797 29515 56831
rect 29457 56791 29515 56797
rect 29549 56831 29607 56837
rect 29549 56797 29561 56831
rect 29595 56797 29607 56831
rect 29549 56791 29607 56797
rect 29641 56831 29699 56837
rect 29641 56797 29653 56831
rect 29687 56797 29699 56831
rect 29822 56828 29828 56840
rect 29783 56800 29828 56828
rect 29641 56791 29699 56797
rect 28074 56760 28080 56772
rect 27816 56732 28080 56760
rect 28074 56720 28080 56732
rect 28132 56720 28138 56772
rect 28534 56720 28540 56772
rect 28592 56760 28598 56772
rect 29549 56760 29577 56791
rect 29822 56788 29828 56800
rect 29880 56788 29886 56840
rect 29932 56760 29960 56868
rect 31113 56865 31125 56899
rect 31159 56896 31171 56899
rect 33704 56896 33732 56936
rect 34790 56924 34796 56936
rect 34848 56924 34854 56976
rect 31159 56868 31892 56896
rect 31159 56865 31171 56868
rect 31113 56859 31171 56865
rect 30929 56831 30987 56837
rect 30929 56797 30941 56831
rect 30975 56797 30987 56831
rect 30929 56791 30987 56797
rect 28592 56732 29960 56760
rect 30944 56760 30972 56791
rect 31018 56788 31024 56840
rect 31076 56828 31082 56840
rect 31205 56831 31263 56837
rect 31076 56800 31121 56828
rect 31076 56788 31082 56800
rect 31205 56797 31217 56831
rect 31251 56828 31263 56831
rect 31754 56828 31760 56840
rect 31251 56800 31760 56828
rect 31251 56797 31263 56800
rect 31205 56791 31263 56797
rect 31754 56788 31760 56800
rect 31812 56788 31818 56840
rect 31864 56828 31892 56868
rect 32324 56868 33456 56896
rect 32324 56837 32352 56868
rect 33428 56840 33456 56868
rect 33612 56868 33732 56896
rect 31938 56831 31996 56837
rect 31938 56828 31950 56831
rect 31864 56800 31950 56828
rect 31938 56797 31950 56800
rect 31984 56828 31996 56831
rect 32309 56831 32367 56837
rect 31984 56800 32260 56828
rect 31984 56797 31996 56800
rect 31938 56791 31996 56797
rect 32232 56772 32260 56800
rect 32309 56797 32321 56831
rect 32355 56797 32367 56831
rect 32309 56791 32367 56797
rect 32401 56831 32459 56837
rect 32401 56797 32413 56831
rect 32447 56822 32459 56831
rect 33410 56828 33416 56840
rect 32447 56797 32536 56822
rect 33371 56800 33416 56828
rect 32401 56794 32536 56797
rect 32401 56791 32459 56794
rect 30944 56732 31984 56760
rect 28592 56720 28598 56732
rect 24121 56695 24179 56701
rect 24121 56661 24133 56695
rect 24167 56692 24179 56695
rect 24486 56692 24492 56704
rect 24167 56664 24492 56692
rect 24167 56661 24179 56664
rect 24121 56655 24179 56661
rect 24486 56652 24492 56664
rect 24544 56652 24550 56704
rect 25038 56652 25044 56704
rect 25096 56692 25102 56704
rect 25133 56695 25191 56701
rect 25133 56692 25145 56695
rect 25096 56664 25145 56692
rect 25096 56652 25102 56664
rect 25133 56661 25145 56664
rect 25179 56661 25191 56695
rect 25133 56655 25191 56661
rect 25317 56695 25375 56701
rect 25317 56661 25329 56695
rect 25363 56692 25375 56695
rect 25498 56692 25504 56704
rect 25363 56664 25504 56692
rect 25363 56661 25375 56664
rect 25317 56655 25375 56661
rect 25498 56652 25504 56664
rect 25556 56652 25562 56704
rect 26878 56692 26884 56704
rect 26839 56664 26884 56692
rect 26878 56652 26884 56664
rect 26936 56652 26942 56704
rect 29089 56695 29147 56701
rect 29089 56661 29101 56695
rect 29135 56692 29147 56695
rect 29454 56692 29460 56704
rect 29135 56664 29460 56692
rect 29135 56661 29147 56664
rect 29089 56655 29147 56661
rect 29454 56652 29460 56664
rect 29512 56652 29518 56704
rect 30006 56652 30012 56704
rect 30064 56692 30070 56704
rect 30745 56695 30803 56701
rect 30745 56692 30757 56695
rect 30064 56664 30757 56692
rect 30064 56652 30070 56664
rect 30745 56661 30757 56664
rect 30791 56661 30803 56695
rect 30745 56655 30803 56661
rect 31754 56652 31760 56704
rect 31812 56692 31818 56704
rect 31956 56701 31984 56732
rect 32214 56720 32220 56772
rect 32272 56720 32278 56772
rect 32508 56760 32536 56794
rect 33410 56788 33416 56800
rect 33468 56788 33474 56840
rect 33505 56831 33563 56837
rect 33505 56797 33517 56831
rect 33551 56828 33563 56831
rect 33612 56828 33640 56868
rect 34330 56856 34336 56908
rect 34388 56896 34394 56908
rect 35161 56899 35219 56905
rect 35161 56896 35173 56899
rect 34388 56868 35173 56896
rect 34388 56856 34394 56868
rect 35161 56865 35173 56868
rect 35207 56865 35219 56899
rect 35161 56859 35219 56865
rect 36173 56899 36231 56905
rect 36173 56865 36185 56899
rect 36219 56896 36231 56899
rect 36219 56868 37412 56896
rect 36219 56865 36231 56868
rect 36173 56859 36231 56865
rect 33551 56800 33640 56828
rect 33689 56831 33747 56837
rect 33551 56797 33563 56800
rect 33505 56791 33563 56797
rect 33689 56797 33701 56831
rect 33735 56797 33747 56831
rect 33689 56791 33747 56797
rect 33704 56760 33732 56791
rect 33778 56788 33784 56840
rect 33836 56828 33842 56840
rect 34422 56828 34428 56840
rect 33836 56800 33881 56828
rect 34383 56800 34428 56828
rect 33836 56788 33842 56800
rect 34422 56788 34428 56800
rect 34480 56788 34486 56840
rect 34606 56828 34612 56840
rect 34567 56800 34612 56828
rect 34606 56788 34612 56800
rect 34664 56788 34670 56840
rect 34701 56831 34759 56837
rect 34701 56797 34713 56831
rect 34747 56797 34759 56831
rect 34701 56791 34759 56797
rect 34440 56760 34468 56788
rect 32508 56732 34468 56760
rect 34716 56760 34744 56791
rect 34882 56788 34888 56840
rect 34940 56828 34946 56840
rect 35989 56831 36047 56837
rect 35989 56828 36001 56831
rect 34940 56800 36001 56828
rect 34940 56788 34946 56800
rect 35989 56797 36001 56800
rect 36035 56797 36047 56831
rect 35989 56791 36047 56797
rect 36541 56831 36599 56837
rect 36541 56797 36553 56831
rect 36587 56797 36599 56831
rect 36541 56791 36599 56797
rect 36817 56831 36875 56837
rect 36817 56797 36829 56831
rect 36863 56828 36875 56831
rect 37274 56828 37280 56840
rect 36863 56800 37280 56828
rect 36863 56797 36875 56800
rect 36817 56791 36875 56797
rect 36446 56760 36452 56772
rect 34716 56732 36452 56760
rect 36446 56720 36452 56732
rect 36504 56720 36510 56772
rect 31941 56695 31999 56701
rect 31812 56664 31857 56692
rect 31812 56652 31818 56664
rect 31941 56661 31953 56695
rect 31987 56692 31999 56695
rect 32030 56692 32036 56704
rect 31987 56664 32036 56692
rect 31987 56661 31999 56664
rect 31941 56655 31999 56661
rect 32030 56652 32036 56664
rect 32088 56652 32094 56704
rect 33226 56692 33232 56704
rect 33187 56664 33232 56692
rect 33226 56652 33232 56664
rect 33284 56652 33290 56704
rect 36078 56692 36084 56704
rect 36039 56664 36084 56692
rect 36078 56652 36084 56664
rect 36136 56652 36142 56704
rect 36556 56692 36584 56791
rect 37274 56788 37280 56800
rect 37332 56788 37338 56840
rect 37384 56828 37412 56868
rect 37461 56831 37519 56837
rect 37461 56828 37473 56831
rect 37384 56800 37473 56828
rect 37461 56797 37473 56800
rect 37507 56828 37519 56831
rect 37568 56828 37596 57004
rect 39758 56964 39764 56976
rect 39040 56936 39764 56964
rect 37826 56856 37832 56908
rect 37884 56896 37890 56908
rect 39040 56905 39068 56936
rect 39758 56924 39764 56936
rect 39816 56924 39822 56976
rect 40402 56924 40408 56976
rect 40460 56924 40466 56976
rect 42889 56967 42947 56973
rect 42889 56964 42901 56967
rect 41708 56936 42901 56964
rect 38657 56899 38715 56905
rect 38657 56896 38669 56899
rect 37884 56868 38669 56896
rect 37884 56856 37890 56868
rect 38657 56865 38669 56868
rect 38703 56865 38715 56899
rect 38657 56859 38715 56865
rect 39025 56899 39083 56905
rect 39025 56865 39037 56899
rect 39071 56865 39083 56899
rect 39025 56859 39083 56865
rect 39117 56899 39175 56905
rect 39117 56865 39129 56899
rect 39163 56896 39175 56899
rect 40420 56896 40448 56924
rect 39163 56868 40448 56896
rect 40773 56899 40831 56905
rect 39163 56865 39175 56868
rect 39117 56859 39175 56865
rect 40773 56865 40785 56899
rect 40819 56896 40831 56899
rect 41708 56896 41736 56936
rect 42889 56933 42901 56936
rect 42935 56964 42947 56967
rect 43806 56964 43812 56976
rect 42935 56936 43812 56964
rect 42935 56933 42947 56936
rect 42889 56927 42947 56933
rect 43806 56924 43812 56936
rect 43864 56924 43870 56976
rect 44284 56973 44312 57004
rect 46014 56992 46020 57044
rect 46072 57032 46078 57044
rect 47581 57035 47639 57041
rect 47581 57032 47593 57035
rect 46072 57004 47593 57032
rect 46072 56992 46078 57004
rect 47581 57001 47593 57004
rect 47627 57001 47639 57035
rect 47581 56995 47639 57001
rect 48774 56992 48780 57044
rect 48832 57032 48838 57044
rect 48869 57035 48927 57041
rect 48869 57032 48881 57035
rect 48832 57004 48881 57032
rect 48832 56992 48838 57004
rect 48869 57001 48881 57004
rect 48915 57001 48927 57035
rect 49694 57032 49700 57044
rect 49655 57004 49700 57032
rect 48869 56995 48927 57001
rect 49694 56992 49700 57004
rect 49752 56992 49758 57044
rect 50154 56992 50160 57044
rect 50212 57032 50218 57044
rect 50341 57035 50399 57041
rect 50341 57032 50353 57035
rect 50212 57004 50353 57032
rect 50212 56992 50218 57004
rect 50341 57001 50353 57004
rect 50387 57001 50399 57035
rect 50341 56995 50399 57001
rect 50614 56992 50620 57044
rect 50672 57032 50678 57044
rect 50985 57035 51043 57041
rect 50985 57032 50997 57035
rect 50672 57004 50997 57032
rect 50672 56992 50678 57004
rect 50985 57001 50997 57004
rect 51031 57001 51043 57035
rect 50985 56995 51043 57001
rect 51534 56992 51540 57044
rect 51592 57032 51598 57044
rect 51629 57035 51687 57041
rect 51629 57032 51641 57035
rect 51592 57004 51641 57032
rect 51592 56992 51598 57004
rect 51629 57001 51641 57004
rect 51675 57001 51687 57035
rect 52454 57032 52460 57044
rect 52415 57004 52460 57032
rect 51629 56995 51687 57001
rect 52454 56992 52460 57004
rect 52512 56992 52518 57044
rect 52914 56992 52920 57044
rect 52972 57032 52978 57044
rect 53101 57035 53159 57041
rect 53101 57032 53113 57035
rect 52972 57004 53113 57032
rect 52972 56992 52978 57004
rect 53101 57001 53113 57004
rect 53147 57001 53159 57035
rect 53101 56995 53159 57001
rect 53374 56992 53380 57044
rect 53432 57032 53438 57044
rect 53745 57035 53803 57041
rect 53745 57032 53757 57035
rect 53432 57004 53757 57032
rect 53432 56992 53438 57004
rect 53745 57001 53757 57004
rect 53791 57001 53803 57035
rect 53745 56995 53803 57001
rect 54294 56992 54300 57044
rect 54352 57032 54358 57044
rect 54389 57035 54447 57041
rect 54389 57032 54401 57035
rect 54352 57004 54401 57032
rect 54352 56992 54358 57004
rect 54389 57001 54401 57004
rect 54435 57001 54447 57035
rect 54389 56995 54447 57001
rect 56134 56992 56140 57044
rect 56192 57032 56198 57044
rect 56229 57035 56287 57041
rect 56229 57032 56241 57035
rect 56192 57004 56241 57032
rect 56192 56992 56198 57004
rect 56229 57001 56241 57004
rect 56275 57001 56287 57035
rect 56229 56995 56287 57001
rect 44269 56967 44327 56973
rect 44269 56933 44281 56967
rect 44315 56933 44327 56967
rect 44269 56927 44327 56933
rect 46934 56924 46940 56976
rect 46992 56964 46998 56976
rect 48225 56967 48283 56973
rect 48225 56964 48237 56967
rect 46992 56936 48237 56964
rect 46992 56924 46998 56936
rect 48225 56933 48237 56936
rect 48271 56933 48283 56967
rect 54110 56964 54116 56976
rect 48225 56927 48283 56933
rect 51046 56936 54116 56964
rect 42981 56899 43039 56905
rect 42981 56896 42993 56899
rect 40819 56868 41736 56896
rect 40819 56865 40831 56868
rect 40773 56859 40831 56865
rect 37507 56800 37596 56828
rect 37737 56831 37795 56837
rect 37507 56797 37519 56800
rect 37461 56791 37519 56797
rect 37737 56797 37749 56831
rect 37783 56797 37795 56831
rect 38838 56828 38844 56840
rect 38799 56800 38844 56828
rect 37737 56791 37795 56797
rect 37292 56760 37320 56788
rect 37752 56760 37780 56791
rect 38838 56788 38844 56800
rect 38896 56788 38902 56840
rect 38930 56788 38936 56840
rect 38988 56828 38994 56840
rect 39761 56831 39819 56837
rect 38988 56800 39033 56828
rect 38988 56788 38994 56800
rect 39761 56797 39773 56831
rect 39807 56828 39819 56831
rect 40126 56828 40132 56840
rect 39807 56800 40132 56828
rect 39807 56797 39819 56800
rect 39761 56791 39819 56797
rect 40126 56788 40132 56800
rect 40184 56788 40190 56840
rect 40218 56788 40224 56840
rect 40276 56828 40282 56840
rect 41708 56837 41736 56868
rect 41800 56868 42993 56896
rect 41800 56840 41828 56868
rect 42981 56865 42993 56868
rect 43027 56896 43039 56899
rect 44174 56896 44180 56908
rect 43027 56868 43576 56896
rect 44135 56868 44180 56896
rect 43027 56865 43039 56868
rect 42981 56859 43039 56865
rect 40346 56831 40404 56837
rect 40346 56828 40358 56831
rect 40276 56800 40358 56828
rect 40276 56788 40282 56800
rect 40346 56797 40358 56800
rect 40392 56797 40404 56831
rect 40346 56791 40404 56797
rect 40865 56831 40923 56837
rect 40865 56797 40877 56831
rect 40911 56797 40923 56831
rect 40865 56791 40923 56797
rect 41693 56831 41751 56837
rect 41693 56797 41705 56831
rect 41739 56797 41751 56831
rect 41693 56791 41751 56797
rect 40880 56760 40908 56791
rect 41782 56788 41788 56840
rect 41840 56828 41846 56840
rect 41969 56831 42027 56837
rect 41840 56800 41933 56828
rect 41840 56788 41846 56800
rect 41969 56797 41981 56831
rect 42015 56797 42027 56831
rect 41969 56791 42027 56797
rect 42061 56831 42119 56837
rect 42061 56797 42073 56831
rect 42107 56828 42119 56831
rect 42521 56831 42579 56837
rect 42521 56828 42533 56831
rect 42107 56800 42533 56828
rect 42107 56797 42119 56800
rect 42061 56791 42119 56797
rect 42521 56797 42533 56800
rect 42567 56797 42579 56831
rect 42702 56828 42708 56840
rect 42663 56800 42708 56828
rect 42521 56791 42579 56797
rect 41984 56760 42012 56791
rect 42702 56788 42708 56800
rect 42760 56788 42766 56840
rect 43438 56828 43444 56840
rect 43399 56800 43444 56828
rect 43438 56788 43444 56800
rect 43496 56788 43502 56840
rect 43548 56828 43576 56868
rect 44174 56856 44180 56868
rect 44232 56856 44238 56908
rect 45002 56896 45008 56908
rect 44915 56868 45008 56896
rect 45002 56856 45008 56868
rect 45060 56896 45066 56908
rect 51046 56896 51074 56936
rect 54110 56924 54116 56936
rect 54168 56924 54174 56976
rect 45060 56868 51074 56896
rect 45060 56856 45066 56868
rect 54754 56856 54760 56908
rect 54812 56896 54818 56908
rect 55217 56899 55275 56905
rect 55217 56896 55229 56899
rect 54812 56868 55229 56896
rect 54812 56856 54818 56868
rect 55217 56865 55229 56868
rect 55263 56865 55275 56899
rect 55217 56859 55275 56865
rect 44082 56828 44088 56840
rect 43548 56800 44088 56828
rect 44082 56788 44088 56800
rect 44140 56788 44146 56840
rect 44361 56831 44419 56837
rect 44361 56797 44373 56831
rect 44407 56797 44419 56831
rect 44726 56828 44732 56840
rect 44687 56800 44732 56828
rect 44361 56791 44419 56797
rect 42150 56760 42156 56772
rect 37292 56732 37780 56760
rect 39500 56732 42156 56760
rect 37645 56695 37703 56701
rect 37645 56692 37657 56695
rect 36556 56664 37657 56692
rect 37645 56661 37657 56664
rect 37691 56692 37703 56695
rect 39500 56692 39528 56732
rect 42150 56720 42156 56732
rect 42208 56760 42214 56772
rect 44376 56760 44404 56791
rect 44726 56788 44732 56800
rect 44784 56788 44790 56840
rect 45646 56828 45652 56840
rect 45607 56800 45652 56828
rect 45646 56788 45652 56800
rect 45704 56788 45710 56840
rect 46106 56828 46112 56840
rect 46067 56800 46112 56828
rect 46106 56788 46112 56800
rect 46164 56788 46170 56840
rect 46934 56828 46940 56840
rect 46895 56800 46940 56828
rect 46934 56788 46940 56800
rect 46992 56788 46998 56840
rect 42208 56732 44404 56760
rect 42208 56720 42214 56732
rect 37691 56664 39528 56692
rect 40221 56695 40279 56701
rect 37691 56661 37703 56664
rect 37645 56655 37703 56661
rect 40221 56661 40233 56695
rect 40267 56692 40279 56695
rect 40310 56692 40316 56704
rect 40267 56664 40316 56692
rect 40267 56661 40279 56664
rect 40221 56655 40279 56661
rect 40310 56652 40316 56664
rect 40368 56652 40374 56704
rect 40405 56695 40463 56701
rect 40405 56661 40417 56695
rect 40451 56692 40463 56695
rect 40586 56692 40592 56704
rect 40451 56664 40592 56692
rect 40451 56661 40463 56664
rect 40405 56655 40463 56661
rect 40586 56652 40592 56664
rect 40644 56652 40650 56704
rect 41322 56652 41328 56704
rect 41380 56692 41386 56704
rect 41509 56695 41567 56701
rect 41509 56692 41521 56695
rect 41380 56664 41521 56692
rect 41380 56652 41386 56664
rect 41509 56661 41521 56664
rect 41555 56661 41567 56695
rect 41509 56655 41567 56661
rect 43162 56652 43168 56704
rect 43220 56692 43226 56704
rect 44744 56692 44772 56788
rect 45462 56692 45468 56704
rect 43220 56664 44772 56692
rect 45423 56664 45468 56692
rect 43220 56652 43226 56664
rect 45462 56652 45468 56664
rect 45520 56652 45526 56704
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 24026 56488 24032 56500
rect 23987 56460 24032 56488
rect 24026 56448 24032 56460
rect 24084 56448 24090 56500
rect 28077 56491 28135 56497
rect 28077 56457 28089 56491
rect 28123 56488 28135 56491
rect 28166 56488 28172 56500
rect 28123 56460 28172 56488
rect 28123 56457 28135 56460
rect 28077 56451 28135 56457
rect 28166 56448 28172 56460
rect 28224 56448 28230 56500
rect 30466 56488 30472 56500
rect 28966 56460 30472 56488
rect 27890 56380 27896 56432
rect 27948 56420 27954 56432
rect 28445 56423 28503 56429
rect 28445 56420 28457 56423
rect 27948 56392 28457 56420
rect 27948 56380 27954 56392
rect 28445 56389 28457 56392
rect 28491 56420 28503 56423
rect 28626 56420 28632 56432
rect 28491 56392 28632 56420
rect 28491 56389 28503 56392
rect 28445 56383 28503 56389
rect 28626 56380 28632 56392
rect 28684 56380 28690 56432
rect 22554 56312 22560 56364
rect 22612 56352 22618 56364
rect 22649 56355 22707 56361
rect 22649 56352 22661 56355
rect 22612 56324 22661 56352
rect 22612 56312 22618 56324
rect 22649 56321 22661 56324
rect 22695 56321 22707 56355
rect 22649 56315 22707 56321
rect 24213 56355 24271 56361
rect 24213 56321 24225 56355
rect 24259 56352 24271 56355
rect 24486 56352 24492 56364
rect 24259 56324 24492 56352
rect 24259 56321 24271 56324
rect 24213 56315 24271 56321
rect 24486 56312 24492 56324
rect 24544 56312 24550 56364
rect 25498 56352 25504 56364
rect 25459 56324 25504 56352
rect 25498 56312 25504 56324
rect 25556 56312 25562 56364
rect 26234 56312 26240 56364
rect 26292 56361 26298 56364
rect 26292 56355 26305 56361
rect 26293 56352 26305 56355
rect 27338 56352 27344 56364
rect 26293 56324 26337 56352
rect 27299 56324 27344 56352
rect 26293 56321 26305 56324
rect 26292 56315 26305 56321
rect 26292 56312 26298 56315
rect 27338 56312 27344 56324
rect 27396 56312 27402 56364
rect 28258 56352 28264 56364
rect 28219 56324 28264 56352
rect 28258 56312 28264 56324
rect 28316 56312 28322 56364
rect 23569 56287 23627 56293
rect 23569 56253 23581 56287
rect 23615 56284 23627 56287
rect 23658 56284 23664 56296
rect 23615 56256 23664 56284
rect 23615 56253 23627 56256
rect 23569 56247 23627 56253
rect 23658 56244 23664 56256
rect 23716 56284 23722 56296
rect 24397 56287 24455 56293
rect 24397 56284 24409 56287
rect 23716 56256 24409 56284
rect 23716 56244 23722 56256
rect 24397 56253 24409 56256
rect 24443 56284 24455 56287
rect 25130 56284 25136 56296
rect 24443 56256 25136 56284
rect 24443 56253 24455 56256
rect 24397 56247 24455 56253
rect 25130 56244 25136 56256
rect 25188 56284 25194 56296
rect 25317 56287 25375 56293
rect 25317 56284 25329 56287
rect 25188 56256 25329 56284
rect 25188 56244 25194 56256
rect 25317 56253 25329 56256
rect 25363 56284 25375 56287
rect 26513 56287 26571 56293
rect 26513 56284 26525 56287
rect 25363 56256 26525 56284
rect 25363 56253 25375 56256
rect 25317 56247 25375 56253
rect 26513 56253 26525 56256
rect 26559 56284 26571 56287
rect 27525 56287 27583 56293
rect 27525 56284 27537 56287
rect 26559 56256 27537 56284
rect 26559 56253 26571 56256
rect 26513 56247 26571 56253
rect 27525 56253 27537 56256
rect 27571 56284 27583 56287
rect 27706 56284 27712 56296
rect 27571 56256 27712 56284
rect 27571 56253 27583 56256
rect 27525 56247 27583 56253
rect 27706 56244 27712 56256
rect 27764 56244 27770 56296
rect 27982 56244 27988 56296
rect 28040 56284 28046 56296
rect 28966 56284 28994 56460
rect 30466 56448 30472 56460
rect 30524 56448 30530 56500
rect 31757 56491 31815 56497
rect 31757 56457 31769 56491
rect 31803 56488 31815 56491
rect 31846 56488 31852 56500
rect 31803 56460 31852 56488
rect 31803 56457 31815 56460
rect 31757 56451 31815 56457
rect 31846 56448 31852 56460
rect 31904 56448 31910 56500
rect 32674 56488 32680 56500
rect 32635 56460 32680 56488
rect 32674 56448 32680 56460
rect 32732 56448 32738 56500
rect 34514 56488 34520 56500
rect 33888 56460 34520 56488
rect 30742 56420 30748 56432
rect 29104 56392 30748 56420
rect 29104 56352 29132 56392
rect 30742 56380 30748 56392
rect 30800 56380 30806 56432
rect 33888 56429 33916 56460
rect 34514 56448 34520 56460
rect 34572 56488 34578 56500
rect 34790 56488 34796 56500
rect 34572 56460 34796 56488
rect 34572 56448 34578 56460
rect 34790 56448 34796 56460
rect 34848 56448 34854 56500
rect 35526 56488 35532 56500
rect 35487 56460 35532 56488
rect 35526 56448 35532 56460
rect 35584 56448 35590 56500
rect 36170 56448 36176 56500
rect 36228 56488 36234 56500
rect 36357 56491 36415 56497
rect 36357 56488 36369 56491
rect 36228 56460 36369 56488
rect 36228 56448 36234 56460
rect 36357 56457 36369 56460
rect 36403 56457 36415 56491
rect 37274 56488 37280 56500
rect 37235 56460 37280 56488
rect 36357 56451 36415 56457
rect 37274 56448 37280 56460
rect 37332 56448 37338 56500
rect 42058 56488 42064 56500
rect 41984 56460 42064 56488
rect 33873 56423 33931 56429
rect 32232 56392 33824 56420
rect 32232 56364 32260 56392
rect 29181 56355 29239 56361
rect 29181 56352 29193 56355
rect 29104 56324 29193 56352
rect 29181 56321 29193 56324
rect 29227 56321 29239 56355
rect 29362 56352 29368 56364
rect 29323 56324 29368 56352
rect 29181 56315 29239 56321
rect 29362 56312 29368 56324
rect 29420 56312 29426 56364
rect 29454 56312 29460 56364
rect 29512 56352 29518 56364
rect 29641 56355 29699 56361
rect 29512 56324 29557 56352
rect 29512 56312 29518 56324
rect 29641 56321 29653 56355
rect 29687 56352 29699 56355
rect 29822 56352 29828 56364
rect 29687 56324 29828 56352
rect 29687 56321 29699 56324
rect 29641 56315 29699 56321
rect 28040 56256 28994 56284
rect 29104 56256 29408 56284
rect 28040 56244 28046 56256
rect 23198 56176 23204 56228
rect 23256 56216 23262 56228
rect 29104 56216 29132 56256
rect 29270 56216 29276 56228
rect 23256 56188 29132 56216
rect 29231 56188 29276 56216
rect 23256 56176 23262 56188
rect 29270 56176 29276 56188
rect 29328 56176 29334 56228
rect 29380 56216 29408 56256
rect 29748 56216 29776 56324
rect 29822 56312 29828 56324
rect 29880 56312 29886 56364
rect 30190 56312 30196 56364
rect 30248 56352 30254 56364
rect 30285 56355 30343 56361
rect 30285 56352 30297 56355
rect 30248 56324 30297 56352
rect 30248 56312 30254 56324
rect 30285 56321 30297 56324
rect 30331 56321 30343 56355
rect 30285 56315 30343 56321
rect 30834 56312 30840 56364
rect 30892 56352 30898 56364
rect 30929 56355 30987 56361
rect 30929 56352 30941 56355
rect 30892 56324 30941 56352
rect 30892 56312 30898 56324
rect 30929 56321 30941 56324
rect 30975 56321 30987 56355
rect 30929 56315 30987 56321
rect 31754 56312 31760 56364
rect 31812 56352 31818 56364
rect 31941 56355 31999 56361
rect 31941 56352 31953 56355
rect 31812 56324 31953 56352
rect 31812 56312 31818 56324
rect 31941 56321 31953 56324
rect 31987 56321 31999 56355
rect 32214 56352 32220 56364
rect 32127 56324 32220 56352
rect 31941 56315 31999 56321
rect 32214 56312 32220 56324
rect 32272 56312 32278 56364
rect 32861 56355 32919 56361
rect 32861 56321 32873 56355
rect 32907 56352 32919 56355
rect 33226 56352 33232 56364
rect 32907 56324 33232 56352
rect 32907 56321 32919 56324
rect 32861 56315 32919 56321
rect 33226 56312 33232 56324
rect 33284 56312 33290 56364
rect 30466 56284 30472 56296
rect 30379 56256 30472 56284
rect 30466 56244 30472 56256
rect 30524 56244 30530 56296
rect 33134 56284 33140 56296
rect 33095 56256 33140 56284
rect 33134 56244 33140 56256
rect 33192 56244 33198 56296
rect 29380 56188 29776 56216
rect 30484 56216 30512 56244
rect 33686 56216 33692 56228
rect 30484 56188 33692 56216
rect 33686 56176 33692 56188
rect 33744 56176 33750 56228
rect 25682 56148 25688 56160
rect 25643 56120 25688 56148
rect 25682 56108 25688 56120
rect 25740 56108 25746 56160
rect 27154 56148 27160 56160
rect 27115 56120 27160 56148
rect 27154 56108 27160 56120
rect 27212 56108 27218 56160
rect 28994 56148 29000 56160
rect 28955 56120 29000 56148
rect 28994 56108 29000 56120
rect 29052 56108 29058 56160
rect 30098 56148 30104 56160
rect 30059 56120 30104 56148
rect 30098 56108 30104 56120
rect 30156 56108 30162 56160
rect 31846 56108 31852 56160
rect 31904 56148 31910 56160
rect 32030 56148 32036 56160
rect 31904 56120 32036 56148
rect 31904 56108 31910 56120
rect 32030 56108 32036 56120
rect 32088 56148 32094 56160
rect 32125 56151 32183 56157
rect 32125 56148 32137 56151
rect 32088 56120 32137 56148
rect 32088 56108 32094 56120
rect 32125 56117 32137 56120
rect 32171 56117 32183 56151
rect 33042 56148 33048 56160
rect 33003 56120 33048 56148
rect 32125 56111 32183 56117
rect 33042 56108 33048 56120
rect 33100 56108 33106 56160
rect 33796 56157 33824 56392
rect 33873 56389 33885 56423
rect 33919 56389 33931 56423
rect 34698 56420 34704 56432
rect 34659 56392 34704 56420
rect 33873 56383 33931 56389
rect 34698 56380 34704 56392
rect 34756 56380 34762 56432
rect 34882 56380 34888 56432
rect 34940 56420 34946 56432
rect 36725 56423 36783 56429
rect 36725 56420 36737 56423
rect 34940 56392 35296 56420
rect 34940 56380 34946 56392
rect 34517 56355 34575 56361
rect 34517 56321 34529 56355
rect 34563 56352 34575 56355
rect 34606 56352 34612 56364
rect 34563 56324 34612 56352
rect 34563 56321 34575 56324
rect 34517 56315 34575 56321
rect 34606 56312 34612 56324
rect 34664 56312 34670 56364
rect 35268 56361 35296 56392
rect 35728 56392 36737 56420
rect 34793 56355 34851 56361
rect 34793 56321 34805 56355
rect 34839 56352 34851 56355
rect 35253 56355 35311 56361
rect 34839 56324 35112 56352
rect 34839 56321 34851 56324
rect 34793 56315 34851 56321
rect 33781 56151 33839 56157
rect 33781 56117 33793 56151
rect 33827 56148 33839 56151
rect 33870 56148 33876 56160
rect 33827 56120 33876 56148
rect 33827 56117 33839 56120
rect 33781 56111 33839 56117
rect 33870 56108 33876 56120
rect 33928 56108 33934 56160
rect 33962 56108 33968 56160
rect 34020 56148 34026 56160
rect 34517 56151 34575 56157
rect 34517 56148 34529 56151
rect 34020 56120 34529 56148
rect 34020 56108 34026 56120
rect 34517 56117 34529 56120
rect 34563 56117 34575 56151
rect 35084 56148 35112 56324
rect 35253 56321 35265 56355
rect 35299 56352 35311 56355
rect 35526 56352 35532 56364
rect 35299 56324 35532 56352
rect 35299 56321 35311 56324
rect 35253 56315 35311 56321
rect 35526 56312 35532 56324
rect 35584 56312 35590 56364
rect 35728 56361 35756 56392
rect 36725 56389 36737 56392
rect 36771 56420 36783 56423
rect 37826 56420 37832 56432
rect 36771 56392 37832 56420
rect 36771 56389 36783 56392
rect 36725 56383 36783 56389
rect 37826 56380 37832 56392
rect 37884 56380 37890 56432
rect 40405 56423 40463 56429
rect 40405 56389 40417 56423
rect 40451 56420 40463 56423
rect 40770 56420 40776 56432
rect 40451 56392 40776 56420
rect 40451 56389 40463 56392
rect 40405 56383 40463 56389
rect 40770 56380 40776 56392
rect 40828 56380 40834 56432
rect 35621 56355 35679 56361
rect 35621 56321 35633 56355
rect 35667 56321 35679 56355
rect 35621 56315 35679 56321
rect 35713 56355 35771 56361
rect 35713 56321 35725 56355
rect 35759 56321 35771 56355
rect 35713 56315 35771 56321
rect 36541 56355 36599 56361
rect 36541 56321 36553 56355
rect 36587 56321 36599 56355
rect 37642 56352 37648 56364
rect 37603 56324 37648 56352
rect 36541 56315 36599 56321
rect 35636 56216 35664 56315
rect 36556 56216 36584 56315
rect 37642 56312 37648 56324
rect 37700 56312 37706 56364
rect 38838 56312 38844 56364
rect 38896 56352 38902 56364
rect 39206 56352 39212 56364
rect 38896 56324 39212 56352
rect 38896 56312 38902 56324
rect 39206 56312 39212 56324
rect 39264 56312 39270 56364
rect 39301 56355 39359 56361
rect 39301 56321 39313 56355
rect 39347 56321 39359 56355
rect 39301 56315 39359 56321
rect 39485 56355 39543 56361
rect 39485 56321 39497 56355
rect 39531 56352 39543 56355
rect 39758 56352 39764 56364
rect 39531 56324 39764 56352
rect 39531 56321 39543 56324
rect 39485 56315 39543 56321
rect 37737 56287 37795 56293
rect 37737 56253 37749 56287
rect 37783 56284 37795 56287
rect 38289 56287 38347 56293
rect 38289 56284 38301 56287
rect 37783 56256 38301 56284
rect 37783 56253 37795 56256
rect 37737 56247 37795 56253
rect 38289 56253 38301 56256
rect 38335 56253 38347 56287
rect 38289 56247 38347 56253
rect 38562 56244 38568 56296
rect 38620 56284 38626 56296
rect 38749 56287 38807 56293
rect 38749 56284 38761 56287
rect 38620 56256 38761 56284
rect 38620 56244 38626 56256
rect 38749 56253 38761 56256
rect 38795 56253 38807 56287
rect 38749 56247 38807 56253
rect 35636 56188 36584 56216
rect 36170 56148 36176 56160
rect 35084 56120 36176 56148
rect 34517 56111 34575 56117
rect 36170 56108 36176 56120
rect 36228 56108 36234 56160
rect 36556 56148 36584 56188
rect 38102 56176 38108 56228
rect 38160 56216 38166 56228
rect 38381 56219 38439 56225
rect 38381 56216 38393 56219
rect 38160 56188 38393 56216
rect 38160 56176 38166 56188
rect 38381 56185 38393 56188
rect 38427 56216 38439 56219
rect 38930 56216 38936 56228
rect 38427 56188 38936 56216
rect 38427 56185 38439 56188
rect 38381 56179 38439 56185
rect 38930 56176 38936 56188
rect 38988 56216 38994 56228
rect 39316 56216 39344 56315
rect 39758 56312 39764 56324
rect 39816 56312 39822 56364
rect 40126 56312 40132 56364
rect 40184 56361 40190 56364
rect 40184 56355 40233 56361
rect 40184 56321 40187 56355
rect 40221 56321 40233 56355
rect 40184 56315 40233 56321
rect 40313 56355 40371 56361
rect 40313 56321 40325 56355
rect 40359 56321 40371 56355
rect 40313 56315 40371 56321
rect 40497 56355 40555 56361
rect 40497 56321 40509 56355
rect 40543 56352 40555 56355
rect 40954 56352 40960 56364
rect 40543 56324 40960 56352
rect 40543 56321 40555 56324
rect 40497 56315 40555 56321
rect 40184 56312 40190 56315
rect 40034 56284 40040 56296
rect 39995 56256 40040 56284
rect 40034 56244 40040 56256
rect 40092 56244 40098 56296
rect 40328 56284 40356 56315
rect 40954 56312 40960 56324
rect 41012 56312 41018 56364
rect 41322 56312 41328 56364
rect 41380 56361 41386 56364
rect 41380 56355 41443 56361
rect 41380 56321 41397 56355
rect 41431 56352 41443 56355
rect 41509 56355 41567 56361
rect 41431 56321 41460 56352
rect 41380 56314 41460 56321
rect 41509 56321 41521 56355
rect 41555 56352 41567 56355
rect 41984 56352 42012 56460
rect 42058 56448 42064 56460
rect 42116 56448 42122 56500
rect 48314 56448 48320 56500
rect 48372 56488 48378 56500
rect 49237 56491 49295 56497
rect 49237 56488 49249 56491
rect 48372 56460 49249 56488
rect 48372 56448 48378 56460
rect 49237 56457 49249 56460
rect 49283 56457 49295 56491
rect 49237 56451 49295 56457
rect 49786 56448 49792 56500
rect 49844 56488 49850 56500
rect 51077 56491 51135 56497
rect 51077 56488 51089 56491
rect 49844 56460 51089 56488
rect 49844 56448 49850 56460
rect 51077 56457 51089 56460
rect 51123 56457 51135 56491
rect 51626 56488 51632 56500
rect 51587 56460 51632 56488
rect 51077 56451 51135 56457
rect 51626 56448 51632 56460
rect 51684 56448 51690 56500
rect 52457 56491 52515 56497
rect 52457 56457 52469 56491
rect 52503 56488 52515 56491
rect 52546 56488 52552 56500
rect 52503 56460 52552 56488
rect 52503 56457 52515 56460
rect 52457 56451 52515 56457
rect 52546 56448 52552 56460
rect 52604 56448 52610 56500
rect 53834 56488 53840 56500
rect 53795 56460 53840 56488
rect 53834 56448 53840 56460
rect 53892 56448 53898 56500
rect 55214 56448 55220 56500
rect 55272 56488 55278 56500
rect 55272 56460 55317 56488
rect 55272 56448 55278 56460
rect 44082 56380 44088 56432
rect 44140 56420 44146 56432
rect 45738 56420 45744 56432
rect 44140 56392 45744 56420
rect 44140 56380 44146 56392
rect 45738 56380 45744 56392
rect 45796 56380 45802 56432
rect 42150 56352 42156 56364
rect 41555 56324 42012 56352
rect 42111 56324 42156 56352
rect 41555 56321 41567 56324
rect 41509 56315 41567 56321
rect 41380 56312 41386 56314
rect 42150 56312 42156 56324
rect 42208 56312 42214 56364
rect 42245 56355 42303 56361
rect 42245 56321 42257 56355
rect 42291 56352 42303 56355
rect 43162 56352 43168 56364
rect 42291 56324 42932 56352
rect 43123 56324 43168 56352
rect 42291 56321 42303 56324
rect 42245 56315 42303 56321
rect 40402 56284 40408 56296
rect 40315 56256 40408 56284
rect 40402 56244 40408 56256
rect 40460 56284 40466 56296
rect 41601 56287 41659 56293
rect 41601 56284 41613 56287
rect 40460 56256 41613 56284
rect 40460 56244 40466 56256
rect 41601 56253 41613 56256
rect 41647 56284 41659 56287
rect 42260 56284 42288 56315
rect 41647 56256 42288 56284
rect 41647 56253 41659 56256
rect 41601 56247 41659 56253
rect 40678 56216 40684 56228
rect 38988 56188 39344 56216
rect 40639 56188 40684 56216
rect 38988 56176 38994 56188
rect 40678 56176 40684 56188
rect 40736 56176 40742 56228
rect 42794 56216 42800 56228
rect 42755 56188 42800 56216
rect 42794 56176 42800 56188
rect 42852 56176 42858 56228
rect 42904 56216 42932 56324
rect 43162 56312 43168 56324
rect 43220 56312 43226 56364
rect 43714 56312 43720 56364
rect 43772 56352 43778 56364
rect 43772 56324 43944 56352
rect 43772 56312 43778 56324
rect 42978 56244 42984 56296
rect 43036 56284 43042 56296
rect 43073 56287 43131 56293
rect 43073 56284 43085 56287
rect 43036 56256 43085 56284
rect 43036 56244 43042 56256
rect 43073 56253 43085 56256
rect 43119 56284 43131 56287
rect 43809 56287 43867 56293
rect 43809 56284 43821 56287
rect 43119 56256 43821 56284
rect 43119 56253 43131 56256
rect 43073 56247 43131 56253
rect 43809 56253 43821 56256
rect 43855 56253 43867 56287
rect 43916 56284 43944 56324
rect 43990 56312 43996 56364
rect 44048 56352 44054 56364
rect 44269 56355 44327 56361
rect 44048 56324 44093 56352
rect 44048 56312 44054 56324
rect 44269 56321 44281 56355
rect 44315 56352 44327 56355
rect 44358 56352 44364 56364
rect 44315 56324 44364 56352
rect 44315 56321 44327 56324
rect 44269 56315 44327 56321
rect 44358 56312 44364 56324
rect 44416 56312 44422 56364
rect 44818 56352 44824 56364
rect 44779 56324 44824 56352
rect 44818 56312 44824 56324
rect 44876 56312 44882 56364
rect 45094 56312 45100 56364
rect 45152 56352 45158 56364
rect 46845 56355 46903 56361
rect 46845 56352 46857 56355
rect 45152 56324 46857 56352
rect 45152 56312 45158 56324
rect 46845 56321 46857 56324
rect 46891 56321 46903 56355
rect 46845 56315 46903 56321
rect 47394 56312 47400 56364
rect 47452 56352 47458 56364
rect 47489 56355 47547 56361
rect 47489 56352 47501 56355
rect 47452 56324 47501 56352
rect 47452 56312 47458 56324
rect 47489 56321 47501 56324
rect 47535 56321 47547 56355
rect 47489 56315 47547 56321
rect 47854 56312 47860 56364
rect 47912 56352 47918 56364
rect 48317 56355 48375 56361
rect 48317 56352 48329 56355
rect 47912 56324 48329 56352
rect 47912 56312 47918 56324
rect 48317 56321 48329 56324
rect 48363 56321 48375 56355
rect 48317 56315 48375 56321
rect 45554 56284 45560 56296
rect 43916 56256 45048 56284
rect 45515 56256 45560 56284
rect 43809 56247 43867 56253
rect 43714 56216 43720 56228
rect 42904 56188 43720 56216
rect 43714 56176 43720 56188
rect 43772 56176 43778 56228
rect 44082 56216 44088 56228
rect 44043 56188 44088 56216
rect 44082 56176 44088 56188
rect 44140 56176 44146 56228
rect 44174 56176 44180 56228
rect 44232 56216 44238 56228
rect 45020 56216 45048 56256
rect 45554 56244 45560 56256
rect 45612 56244 45618 56296
rect 46201 56219 46259 56225
rect 46201 56216 46213 56219
rect 44232 56188 44956 56216
rect 45020 56188 46213 56216
rect 44232 56176 44238 56188
rect 39485 56151 39543 56157
rect 39485 56148 39497 56151
rect 36556 56120 39497 56148
rect 39485 56117 39497 56120
rect 39531 56117 39543 56151
rect 41138 56148 41144 56160
rect 41099 56120 41144 56148
rect 39485 56111 39543 56117
rect 41138 56108 41144 56120
rect 41196 56108 41202 56160
rect 41598 56108 41604 56160
rect 41656 56148 41662 56160
rect 42702 56148 42708 56160
rect 41656 56120 42708 56148
rect 41656 56108 41662 56120
rect 42702 56108 42708 56120
rect 42760 56148 42766 56160
rect 44818 56148 44824 56160
rect 42760 56120 44824 56148
rect 42760 56108 42766 56120
rect 44818 56108 44824 56120
rect 44876 56108 44882 56160
rect 44928 56148 44956 56188
rect 46201 56185 46213 56188
rect 46247 56185 46259 56219
rect 46201 56179 46259 56185
rect 47210 56148 47216 56160
rect 44928 56120 47216 56148
rect 47210 56108 47216 56120
rect 47268 56108 47274 56160
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 23109 55947 23167 55953
rect 23109 55913 23121 55947
rect 23155 55944 23167 55947
rect 23658 55944 23664 55956
rect 23155 55916 23664 55944
rect 23155 55913 23167 55916
rect 23109 55907 23167 55913
rect 23658 55904 23664 55916
rect 23716 55904 23722 55956
rect 23750 55904 23756 55956
rect 23808 55944 23814 55956
rect 24121 55947 24179 55953
rect 24121 55944 24133 55947
rect 23808 55916 24133 55944
rect 23808 55904 23814 55916
rect 24121 55913 24133 55916
rect 24167 55913 24179 55947
rect 24121 55907 24179 55913
rect 25774 55904 25780 55956
rect 25832 55944 25838 55956
rect 26053 55947 26111 55953
rect 26053 55944 26065 55947
rect 25832 55916 26065 55944
rect 25832 55904 25838 55916
rect 26053 55913 26065 55916
rect 26099 55913 26111 55947
rect 28994 55944 29000 55956
rect 26053 55907 26111 55913
rect 26160 55916 29000 55944
rect 17402 55836 17408 55888
rect 17460 55876 17466 55888
rect 26160 55876 26188 55916
rect 28994 55904 29000 55916
rect 29052 55904 29058 55956
rect 30190 55904 30196 55956
rect 30248 55944 30254 55956
rect 34241 55947 34299 55953
rect 34241 55944 34253 55947
rect 30248 55916 34253 55944
rect 30248 55904 30254 55916
rect 34241 55913 34253 55916
rect 34287 55913 34299 55947
rect 34241 55907 34299 55913
rect 34422 55904 34428 55956
rect 34480 55944 34486 55956
rect 35253 55947 35311 55953
rect 35253 55944 35265 55947
rect 34480 55916 35265 55944
rect 34480 55904 34486 55916
rect 35253 55913 35265 55916
rect 35299 55913 35311 55947
rect 39206 55944 39212 55956
rect 35253 55907 35311 55913
rect 36280 55916 39068 55944
rect 39167 55916 39212 55944
rect 17460 55848 26188 55876
rect 27065 55879 27123 55885
rect 17460 55836 17466 55848
rect 27065 55845 27077 55879
rect 27111 55876 27123 55879
rect 28258 55876 28264 55888
rect 27111 55848 28264 55876
rect 27111 55845 27123 55848
rect 27065 55839 27123 55845
rect 28258 55836 28264 55848
rect 28316 55836 28322 55888
rect 28626 55876 28632 55888
rect 28587 55848 28632 55876
rect 28626 55836 28632 55848
rect 28684 55836 28690 55888
rect 33962 55876 33968 55888
rect 29012 55848 33968 55876
rect 27154 55808 27160 55820
rect 25240 55780 27160 55808
rect 24302 55740 24308 55752
rect 24263 55712 24308 55740
rect 24302 55700 24308 55712
rect 24360 55700 24366 55752
rect 25240 55749 25268 55780
rect 27154 55768 27160 55780
rect 27212 55768 27218 55820
rect 27522 55768 27528 55820
rect 27580 55808 27586 55820
rect 29012 55817 29040 55848
rect 33962 55836 33968 55848
rect 34020 55836 34026 55888
rect 34054 55836 34060 55888
rect 34112 55876 34118 55888
rect 35986 55876 35992 55888
rect 34112 55848 35992 55876
rect 34112 55836 34118 55848
rect 35986 55836 35992 55848
rect 36044 55836 36050 55888
rect 28997 55811 29055 55817
rect 28997 55808 29009 55811
rect 27580 55780 29009 55808
rect 27580 55768 27586 55780
rect 28997 55777 29009 55780
rect 29043 55777 29055 55811
rect 28997 55771 29055 55777
rect 29089 55811 29147 55817
rect 29089 55777 29101 55811
rect 29135 55808 29147 55811
rect 29178 55808 29184 55820
rect 29135 55780 29184 55808
rect 29135 55777 29147 55780
rect 29089 55771 29147 55777
rect 29178 55768 29184 55780
rect 29236 55808 29242 55820
rect 30374 55808 30380 55820
rect 29236 55780 30380 55808
rect 29236 55768 29242 55780
rect 30374 55768 30380 55780
rect 30432 55808 30438 55820
rect 31018 55808 31024 55820
rect 30432 55780 31024 55808
rect 30432 55768 30438 55780
rect 31018 55768 31024 55780
rect 31076 55808 31082 55820
rect 33505 55811 33563 55817
rect 33505 55808 33517 55811
rect 31076 55780 31156 55808
rect 31076 55768 31082 55780
rect 25225 55743 25283 55749
rect 25225 55709 25237 55743
rect 25271 55709 25283 55743
rect 25866 55740 25872 55752
rect 25827 55712 25872 55740
rect 25225 55703 25283 55709
rect 25866 55700 25872 55712
rect 25924 55700 25930 55752
rect 26789 55743 26847 55749
rect 26789 55709 26801 55743
rect 26835 55740 26847 55743
rect 28810 55740 28816 55752
rect 26835 55712 27660 55740
rect 26835 55709 26847 55712
rect 26789 55703 26847 55709
rect 27065 55675 27123 55681
rect 27065 55641 27077 55675
rect 27111 55672 27123 55675
rect 27522 55672 27528 55684
rect 27111 55644 27528 55672
rect 27111 55641 27123 55644
rect 27065 55635 27123 55641
rect 27522 55632 27528 55644
rect 27580 55632 27586 55684
rect 27632 55672 27660 55712
rect 27816 55712 28816 55740
rect 27816 55672 27844 55712
rect 28810 55700 28816 55712
rect 28868 55700 28874 55752
rect 28902 55700 28908 55752
rect 28960 55740 28966 55752
rect 29638 55740 29644 55752
rect 28960 55712 29005 55740
rect 29599 55712 29644 55740
rect 28960 55700 28966 55712
rect 29638 55700 29644 55712
rect 29696 55700 29702 55752
rect 30282 55700 30288 55752
rect 30340 55740 30346 55752
rect 31128 55749 31156 55780
rect 31726 55780 33517 55808
rect 30837 55743 30895 55749
rect 30837 55740 30849 55743
rect 30340 55712 30849 55740
rect 30340 55700 30346 55712
rect 30837 55709 30849 55712
rect 30883 55709 30895 55743
rect 30837 55703 30895 55709
rect 31113 55743 31171 55749
rect 31113 55709 31125 55743
rect 31159 55709 31171 55743
rect 31113 55703 31171 55709
rect 31297 55743 31355 55749
rect 31297 55709 31309 55743
rect 31343 55740 31355 55743
rect 31726 55740 31754 55780
rect 33505 55777 33517 55780
rect 33551 55777 33563 55811
rect 33505 55771 33563 55777
rect 34606 55768 34612 55820
rect 34664 55808 34670 55820
rect 36078 55808 36084 55820
rect 34664 55780 34709 55808
rect 35360 55780 36084 55808
rect 34664 55768 34670 55780
rect 32122 55740 32128 55752
rect 31343 55712 31754 55740
rect 32083 55712 32128 55740
rect 31343 55709 31355 55712
rect 31297 55703 31355 55709
rect 32122 55700 32128 55712
rect 32180 55700 32186 55752
rect 32398 55740 32404 55752
rect 32359 55712 32404 55740
rect 32398 55700 32404 55712
rect 32456 55740 32462 55752
rect 33137 55743 33195 55749
rect 33137 55740 33149 55743
rect 32456 55712 33149 55740
rect 32456 55700 32462 55712
rect 33137 55709 33149 55712
rect 33183 55709 33195 55743
rect 33137 55703 33195 55709
rect 33321 55743 33379 55749
rect 33321 55709 33333 55743
rect 33367 55740 33379 55743
rect 33410 55740 33416 55752
rect 33367 55712 33416 55740
rect 33367 55709 33379 55712
rect 33321 55703 33379 55709
rect 27982 55672 27988 55684
rect 27632 55644 27844 55672
rect 27943 55644 27988 55672
rect 27982 55632 27988 55644
rect 28040 55632 28046 55684
rect 28169 55675 28227 55681
rect 28169 55641 28181 55675
rect 28215 55672 28227 55675
rect 30190 55672 30196 55684
rect 28215 55644 30196 55672
rect 28215 55641 28227 55644
rect 28169 55635 28227 55641
rect 30190 55632 30196 55644
rect 30248 55632 30254 55684
rect 30926 55632 30932 55684
rect 30984 55681 30990 55684
rect 30984 55675 31033 55681
rect 30984 55641 30987 55675
rect 31021 55641 31033 55675
rect 30984 55635 31033 55641
rect 31205 55675 31263 55681
rect 31205 55641 31217 55675
rect 31251 55672 31263 55675
rect 31941 55675 31999 55681
rect 31941 55672 31953 55675
rect 31251 55644 31953 55672
rect 31251 55641 31263 55644
rect 31205 55635 31263 55641
rect 31941 55641 31953 55644
rect 31987 55641 31999 55675
rect 33336 55672 33364 55703
rect 33410 55700 33416 55712
rect 33468 55700 33474 55752
rect 34439 55743 34497 55749
rect 34439 55709 34451 55743
rect 34485 55740 34497 55743
rect 34698 55740 34704 55752
rect 34485 55712 34704 55740
rect 34485 55709 34497 55712
rect 34439 55703 34497 55709
rect 34698 55700 34704 55712
rect 34756 55700 34762 55752
rect 35360 55749 35388 55780
rect 36078 55768 36084 55780
rect 36136 55808 36142 55820
rect 36280 55808 36308 55916
rect 38010 55876 38016 55888
rect 36832 55848 38016 55876
rect 36832 55817 36860 55848
rect 38010 55836 38016 55848
rect 38068 55836 38074 55888
rect 38286 55836 38292 55888
rect 38344 55876 38350 55888
rect 39040 55876 39068 55916
rect 39206 55904 39212 55916
rect 39264 55904 39270 55956
rect 40494 55944 40500 55956
rect 40455 55916 40500 55944
rect 40494 55904 40500 55916
rect 40552 55904 40558 55956
rect 40954 55904 40960 55956
rect 41012 55944 41018 55956
rect 43625 55947 43683 55953
rect 43625 55944 43637 55947
rect 41012 55916 43637 55944
rect 41012 55904 41018 55916
rect 43625 55913 43637 55916
rect 43671 55913 43683 55947
rect 44358 55944 44364 55956
rect 44319 55916 44364 55944
rect 43625 55907 43683 55913
rect 44358 55904 44364 55916
rect 44416 55904 44422 55956
rect 44634 55904 44640 55956
rect 44692 55944 44698 55956
rect 45649 55947 45707 55953
rect 45649 55944 45661 55947
rect 44692 55916 45661 55944
rect 44692 55904 44698 55916
rect 45649 55913 45661 55916
rect 45695 55913 45707 55947
rect 45649 55907 45707 55913
rect 45830 55904 45836 55956
rect 45888 55944 45894 55956
rect 46937 55947 46995 55953
rect 46937 55944 46949 55947
rect 45888 55916 46949 55944
rect 45888 55904 45894 55916
rect 46937 55913 46949 55916
rect 46983 55913 46995 55947
rect 46937 55907 46995 55913
rect 47026 55904 47032 55956
rect 47084 55944 47090 55956
rect 47857 55947 47915 55953
rect 47857 55944 47869 55947
rect 47084 55916 47869 55944
rect 47084 55904 47090 55916
rect 47857 55913 47869 55916
rect 47903 55913 47915 55947
rect 47857 55907 47915 55913
rect 40129 55879 40187 55885
rect 38344 55848 38976 55876
rect 39040 55848 39620 55876
rect 38344 55836 38350 55848
rect 36136 55780 36308 55808
rect 36136 55768 36142 55780
rect 36280 55749 36308 55780
rect 36817 55811 36875 55817
rect 36817 55777 36829 55811
rect 36863 55777 36875 55811
rect 36817 55771 36875 55777
rect 37185 55811 37243 55817
rect 37185 55777 37197 55811
rect 37231 55808 37243 55811
rect 38562 55808 38568 55820
rect 37231 55780 38568 55808
rect 37231 55777 37243 55780
rect 37185 55771 37243 55777
rect 38562 55768 38568 55780
rect 38620 55808 38626 55820
rect 38948 55808 38976 55848
rect 38620 55780 38792 55808
rect 38948 55780 39068 55808
rect 38620 55768 38626 55780
rect 35345 55743 35403 55749
rect 35345 55709 35357 55743
rect 35391 55709 35403 55743
rect 35345 55703 35403 55709
rect 36172 55743 36230 55749
rect 36172 55709 36184 55743
rect 36218 55709 36230 55743
rect 36172 55703 36230 55709
rect 36265 55743 36323 55749
rect 36265 55709 36277 55743
rect 36311 55709 36323 55743
rect 36998 55740 37004 55752
rect 36959 55712 37004 55740
rect 36265 55703 36323 55709
rect 31941 55635 31999 55641
rect 32324 55644 33364 55672
rect 30984 55632 30990 55635
rect 25409 55607 25467 55613
rect 25409 55573 25421 55607
rect 25455 55604 25467 55607
rect 26510 55604 26516 55616
rect 25455 55576 26516 55604
rect 25455 55573 25467 55576
rect 25409 55567 25467 55573
rect 26510 55564 26516 55576
rect 26568 55564 26574 55616
rect 26881 55607 26939 55613
rect 26881 55573 26893 55607
rect 26927 55604 26939 55607
rect 27801 55607 27859 55613
rect 27801 55604 27813 55607
rect 26927 55576 27813 55604
rect 26927 55573 26939 55576
rect 26881 55567 26939 55573
rect 27801 55573 27813 55576
rect 27847 55604 27859 55607
rect 28258 55604 28264 55616
rect 27847 55576 28264 55604
rect 27847 55573 27859 55576
rect 27801 55567 27859 55573
rect 28258 55564 28264 55576
rect 28316 55604 28322 55616
rect 28902 55604 28908 55616
rect 28316 55576 28908 55604
rect 28316 55564 28322 55576
rect 28902 55564 28908 55576
rect 28960 55564 28966 55616
rect 29822 55604 29828 55616
rect 29783 55576 29828 55604
rect 29822 55564 29828 55576
rect 29880 55564 29886 55616
rect 30006 55564 30012 55616
rect 30064 55604 30070 55616
rect 32324 55613 32352 55644
rect 31481 55607 31539 55613
rect 31481 55604 31493 55607
rect 30064 55576 31493 55604
rect 30064 55564 30070 55576
rect 31481 55573 31493 55576
rect 31527 55573 31539 55607
rect 31481 55567 31539 55573
rect 32309 55607 32367 55613
rect 32309 55573 32321 55607
rect 32355 55573 32367 55607
rect 32309 55567 32367 55573
rect 33134 55564 33140 55616
rect 33192 55604 33198 55616
rect 35360 55604 35388 55703
rect 36188 55672 36216 55703
rect 36998 55700 37004 55712
rect 37056 55700 37062 55752
rect 37642 55740 37648 55752
rect 37603 55712 37648 55740
rect 37642 55700 37648 55712
rect 37700 55700 37706 55752
rect 37829 55743 37887 55749
rect 37829 55709 37841 55743
rect 37875 55709 37887 55743
rect 37829 55703 37887 55709
rect 38105 55743 38163 55749
rect 38105 55709 38117 55743
rect 38151 55740 38163 55743
rect 38286 55740 38292 55752
rect 38151 55712 38292 55740
rect 38151 55709 38163 55712
rect 38105 55703 38163 55709
rect 36446 55672 36452 55684
rect 36188 55644 36452 55672
rect 36446 55632 36452 55644
rect 36504 55632 36510 55684
rect 37844 55672 37872 55703
rect 38286 55700 38292 55712
rect 38344 55700 38350 55752
rect 38764 55749 38792 55780
rect 38657 55743 38715 55749
rect 38657 55740 38669 55743
rect 38396 55712 38669 55740
rect 37918 55672 37924 55684
rect 37831 55644 37924 55672
rect 37918 55632 37924 55644
rect 37976 55672 37982 55684
rect 38396 55672 38424 55712
rect 38657 55709 38669 55712
rect 38703 55709 38715 55743
rect 38657 55703 38715 55709
rect 38763 55743 38821 55749
rect 38763 55709 38775 55743
rect 38809 55709 38821 55743
rect 38930 55740 38936 55752
rect 38891 55712 38936 55740
rect 38763 55703 38821 55709
rect 38930 55700 38936 55712
rect 38988 55700 38994 55752
rect 39040 55749 39068 55780
rect 39025 55743 39083 55749
rect 39025 55709 39037 55743
rect 39071 55740 39083 55743
rect 39482 55740 39488 55752
rect 39071 55712 39488 55740
rect 39071 55709 39083 55712
rect 39025 55703 39083 55709
rect 39482 55700 39488 55712
rect 39540 55700 39546 55752
rect 37976 55644 38424 55672
rect 39592 55672 39620 55848
rect 40129 55845 40141 55879
rect 40175 55876 40187 55879
rect 40586 55876 40592 55888
rect 40175 55848 40592 55876
rect 40175 55845 40187 55848
rect 40129 55839 40187 55845
rect 40586 55836 40592 55848
rect 40644 55836 40650 55888
rect 44910 55876 44916 55888
rect 40880 55848 44916 55876
rect 40037 55811 40095 55817
rect 40037 55777 40049 55811
rect 40083 55808 40095 55811
rect 40218 55808 40224 55820
rect 40083 55780 40224 55808
rect 40083 55777 40095 55780
rect 40037 55771 40095 55777
rect 40218 55768 40224 55780
rect 40276 55768 40282 55820
rect 40310 55740 40316 55752
rect 40271 55712 40316 55740
rect 40310 55700 40316 55712
rect 40368 55700 40374 55752
rect 40880 55672 40908 55848
rect 44910 55836 44916 55848
rect 44968 55836 44974 55888
rect 45094 55836 45100 55888
rect 45152 55876 45158 55888
rect 51074 55876 51080 55888
rect 45152 55848 51080 55876
rect 45152 55836 45158 55848
rect 51074 55836 51080 55848
rect 51132 55836 51138 55888
rect 41782 55768 41788 55820
rect 41840 55808 41846 55820
rect 41840 55780 42784 55808
rect 41840 55768 41846 55780
rect 41598 55740 41604 55752
rect 41559 55712 41604 55740
rect 41598 55700 41604 55712
rect 41656 55700 41662 55752
rect 41877 55743 41935 55749
rect 41877 55709 41889 55743
rect 41923 55740 41935 55743
rect 42242 55740 42248 55752
rect 41923 55712 42248 55740
rect 41923 55709 41935 55712
rect 41877 55703 41935 55709
rect 42242 55700 42248 55712
rect 42300 55700 42306 55752
rect 42518 55740 42524 55752
rect 42479 55712 42524 55740
rect 42518 55700 42524 55712
rect 42576 55700 42582 55752
rect 42756 55749 42784 55780
rect 43346 55768 43352 55820
rect 43404 55808 43410 55820
rect 46385 55811 46443 55817
rect 43404 55780 45232 55808
rect 43404 55768 43410 55780
rect 42741 55743 42799 55749
rect 42613 55721 42671 55727
rect 42613 55687 42625 55721
rect 42659 55687 42671 55721
rect 42741 55709 42753 55743
rect 42787 55709 42799 55743
rect 42741 55703 42799 55709
rect 43622 55700 43628 55752
rect 43680 55740 43686 55752
rect 43806 55740 43812 55752
rect 43680 55712 43812 55740
rect 43680 55700 43686 55712
rect 43806 55700 43812 55712
rect 43864 55740 43870 55752
rect 45204 55749 45232 55780
rect 46385 55777 46397 55811
rect 46431 55808 46443 55811
rect 50062 55808 50068 55820
rect 46431 55780 50068 55808
rect 46431 55777 46443 55780
rect 46385 55771 46443 55777
rect 44452 55743 44510 55749
rect 44452 55740 44464 55743
rect 43864 55712 44464 55740
rect 43864 55700 43870 55712
rect 44452 55709 44464 55712
rect 44498 55709 44510 55743
rect 44452 55703 44510 55709
rect 44545 55743 44603 55749
rect 44545 55709 44557 55743
rect 44591 55740 44603 55743
rect 45189 55743 45247 55749
rect 44591 55712 44864 55740
rect 44591 55709 44603 55712
rect 44545 55703 44603 55709
rect 42613 55684 42671 55687
rect 39592 55644 40908 55672
rect 37976 55632 37982 55644
rect 42610 55632 42616 55684
rect 42668 55632 42674 55684
rect 43070 55632 43076 55684
rect 43128 55672 43134 55684
rect 43257 55675 43315 55681
rect 43257 55672 43269 55675
rect 43128 55644 43269 55672
rect 43128 55632 43134 55644
rect 43257 55641 43269 55644
rect 43303 55641 43315 55675
rect 43257 55635 43315 55641
rect 43441 55675 43499 55681
rect 43441 55641 43453 55675
rect 43487 55641 43499 55675
rect 43441 55635 43499 55641
rect 33192 55576 35388 55604
rect 35897 55607 35955 55613
rect 33192 55564 33198 55576
rect 35897 55573 35909 55607
rect 35943 55604 35955 55607
rect 36170 55604 36176 55616
rect 35943 55576 36176 55604
rect 35943 55573 35955 55576
rect 35897 55567 35955 55573
rect 36170 55564 36176 55576
rect 36228 55564 36234 55616
rect 38013 55607 38071 55613
rect 38013 55573 38025 55607
rect 38059 55604 38071 55607
rect 38930 55604 38936 55616
rect 38059 55576 38936 55604
rect 38059 55573 38071 55576
rect 38013 55567 38071 55573
rect 38930 55564 38936 55576
rect 38988 55564 38994 55616
rect 41414 55564 41420 55616
rect 41472 55604 41478 55616
rect 41785 55607 41843 55613
rect 41472 55576 41517 55604
rect 41472 55564 41478 55576
rect 41785 55573 41797 55607
rect 41831 55604 41843 55607
rect 41966 55604 41972 55616
rect 41831 55576 41972 55604
rect 41831 55573 41843 55576
rect 41785 55567 41843 55573
rect 41966 55564 41972 55576
rect 42024 55604 42030 55616
rect 42337 55607 42395 55613
rect 42337 55604 42349 55607
rect 42024 55576 42349 55604
rect 42024 55564 42030 55576
rect 42337 55573 42349 55576
rect 42383 55573 42395 55607
rect 43456 55604 43484 55635
rect 43622 55604 43628 55616
rect 43456 55576 43628 55604
rect 42337 55567 42395 55573
rect 43622 55564 43628 55576
rect 43680 55564 43686 55616
rect 43714 55564 43720 55616
rect 43772 55604 43778 55616
rect 44560 55604 44588 55703
rect 44836 55672 44864 55712
rect 45189 55709 45201 55743
rect 45235 55740 45247 55743
rect 45554 55740 45560 55752
rect 45235 55712 45560 55740
rect 45235 55709 45247 55712
rect 45189 55703 45247 55709
rect 45554 55700 45560 55712
rect 45612 55700 45618 55752
rect 46400 55672 46428 55771
rect 50062 55768 50068 55780
rect 50120 55768 50126 55820
rect 44836 55644 46428 55672
rect 43772 55576 44588 55604
rect 43772 55564 43778 55576
rect 44818 55564 44824 55616
rect 44876 55604 44882 55616
rect 45005 55607 45063 55613
rect 45005 55604 45017 55607
rect 44876 55576 45017 55604
rect 44876 55564 44882 55576
rect 45005 55573 45017 55576
rect 45051 55573 45063 55607
rect 45005 55567 45063 55573
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 25406 55360 25412 55412
rect 25464 55400 25470 55412
rect 25501 55403 25559 55409
rect 25501 55400 25513 55403
rect 25464 55372 25513 55400
rect 25464 55360 25470 55372
rect 25501 55369 25513 55372
rect 25547 55369 25559 55403
rect 25501 55363 25559 55369
rect 27338 55360 27344 55412
rect 27396 55400 27402 55412
rect 30006 55400 30012 55412
rect 27396 55372 30012 55400
rect 27396 55360 27402 55372
rect 30006 55360 30012 55372
rect 30064 55360 30070 55412
rect 30098 55360 30104 55412
rect 30156 55360 30162 55412
rect 30282 55409 30288 55412
rect 30278 55400 30288 55409
rect 30243 55372 30288 55400
rect 30278 55363 30288 55372
rect 30282 55360 30288 55363
rect 30340 55360 30346 55412
rect 30837 55403 30895 55409
rect 30837 55369 30849 55403
rect 30883 55400 30895 55403
rect 30926 55400 30932 55412
rect 30883 55372 30932 55400
rect 30883 55369 30895 55372
rect 30837 55363 30895 55369
rect 30926 55360 30932 55372
rect 30984 55360 30990 55412
rect 34517 55403 34575 55409
rect 34517 55369 34529 55403
rect 34563 55400 34575 55403
rect 34606 55400 34612 55412
rect 34563 55372 34612 55400
rect 34563 55369 34575 55372
rect 34517 55363 34575 55369
rect 34606 55360 34612 55372
rect 34664 55360 34670 55412
rect 35618 55400 35624 55412
rect 34716 55372 35624 55400
rect 27985 55335 28043 55341
rect 27985 55301 27997 55335
rect 28031 55332 28043 55335
rect 30116 55332 30144 55360
rect 28031 55304 30144 55332
rect 30193 55335 30251 55341
rect 28031 55301 28043 55304
rect 27985 55295 28043 55301
rect 25682 55264 25688 55276
rect 25643 55236 25688 55264
rect 25682 55224 25688 55236
rect 25740 55224 25746 55276
rect 26234 55224 26240 55276
rect 26292 55264 26298 55276
rect 27065 55267 27123 55273
rect 27065 55264 27077 55267
rect 26292 55236 27077 55264
rect 26292 55224 26298 55236
rect 27065 55233 27077 55236
rect 27111 55233 27123 55267
rect 27065 55227 27123 55233
rect 29178 55224 29184 55276
rect 29236 55264 29242 55276
rect 29273 55267 29331 55273
rect 29273 55264 29285 55267
rect 29236 55236 29285 55264
rect 29236 55224 29242 55236
rect 29273 55233 29285 55236
rect 29319 55233 29331 55267
rect 29273 55227 29331 55233
rect 23934 55156 23940 55208
rect 23992 55196 23998 55208
rect 24029 55199 24087 55205
rect 24029 55196 24041 55199
rect 23992 55168 24041 55196
rect 23992 55156 23998 55168
rect 24029 55165 24041 55168
rect 24075 55165 24087 55199
rect 24029 55159 24087 55165
rect 25041 55199 25099 55205
rect 25041 55165 25053 55199
rect 25087 55196 25099 55199
rect 25314 55196 25320 55208
rect 25087 55168 25320 55196
rect 25087 55165 25099 55168
rect 25041 55159 25099 55165
rect 25314 55156 25320 55168
rect 25372 55156 25378 55208
rect 26605 55199 26663 55205
rect 26605 55165 26617 55199
rect 26651 55196 26663 55199
rect 27798 55196 27804 55208
rect 26651 55168 27804 55196
rect 26651 55165 26663 55168
rect 26605 55159 26663 55165
rect 27798 55156 27804 55168
rect 27856 55156 27862 55208
rect 28810 55156 28816 55208
rect 28868 55196 28874 55208
rect 29089 55199 29147 55205
rect 29089 55196 29101 55199
rect 28868 55168 29101 55196
rect 28868 55156 28874 55168
rect 29089 55165 29101 55168
rect 29135 55165 29147 55199
rect 29288 55196 29316 55227
rect 29362 55224 29368 55276
rect 29420 55264 29426 55276
rect 29561 55273 29589 55304
rect 30193 55301 30205 55335
rect 30239 55332 30251 55335
rect 30466 55332 30472 55344
rect 30239 55304 30472 55332
rect 30239 55301 30251 55304
rect 30193 55295 30251 55301
rect 30466 55292 30472 55304
rect 30524 55332 30530 55344
rect 31021 55335 31079 55341
rect 31021 55332 31033 55335
rect 30524 55304 31033 55332
rect 30524 55292 30530 55304
rect 31021 55301 31033 55304
rect 31067 55301 31079 55335
rect 31021 55295 31079 55301
rect 32122 55292 32128 55344
rect 32180 55332 32186 55344
rect 34716 55332 34744 55372
rect 35618 55360 35624 55372
rect 35676 55360 35682 55412
rect 37918 55360 37924 55412
rect 37976 55400 37982 55412
rect 38013 55403 38071 55409
rect 38013 55400 38025 55403
rect 37976 55372 38025 55400
rect 37976 55360 37982 55372
rect 38013 55369 38025 55372
rect 38059 55369 38071 55403
rect 38013 55363 38071 55369
rect 41601 55403 41659 55409
rect 41601 55369 41613 55403
rect 41647 55400 41659 55403
rect 41782 55400 41788 55412
rect 41647 55372 41788 55400
rect 41647 55369 41659 55372
rect 41601 55363 41659 55369
rect 41782 55360 41788 55372
rect 41840 55360 41846 55412
rect 42518 55360 42524 55412
rect 42576 55400 42582 55412
rect 44358 55400 44364 55412
rect 42576 55372 44364 55400
rect 42576 55360 42582 55372
rect 32180 55304 34744 55332
rect 32180 55292 32186 55304
rect 29508 55267 29589 55273
rect 29420 55236 29465 55264
rect 29420 55224 29426 55236
rect 29508 55233 29520 55267
rect 29554 55234 29589 55267
rect 29651 55267 29709 55273
rect 29554 55233 29566 55234
rect 29508 55227 29566 55233
rect 29651 55233 29663 55267
rect 29697 55264 29709 55267
rect 30006 55264 30012 55276
rect 29697 55236 30012 55264
rect 29697 55233 29709 55236
rect 29651 55227 29709 55233
rect 30006 55224 30012 55236
rect 30064 55224 30070 55276
rect 30101 55267 30159 55273
rect 30101 55233 30113 55267
rect 30147 55233 30159 55267
rect 30374 55264 30380 55276
rect 30335 55236 30380 55264
rect 30101 55227 30159 55233
rect 30116 55196 30144 55227
rect 30374 55224 30380 55236
rect 30432 55224 30438 55276
rect 31205 55267 31263 55273
rect 31205 55233 31217 55267
rect 31251 55233 31263 55267
rect 31205 55227 31263 55233
rect 31849 55267 31907 55273
rect 31849 55233 31861 55267
rect 31895 55264 31907 55267
rect 32214 55264 32220 55276
rect 31895 55236 32220 55264
rect 31895 55233 31907 55236
rect 31849 55227 31907 55233
rect 30282 55196 30288 55208
rect 29288 55168 30288 55196
rect 29089 55159 29147 55165
rect 30282 55156 30288 55168
rect 30340 55196 30346 55208
rect 31220 55196 31248 55227
rect 32214 55224 32220 55236
rect 32272 55224 32278 55276
rect 32766 55224 32772 55276
rect 32824 55264 32830 55276
rect 32824 55236 33088 55264
rect 32824 55224 32830 55236
rect 30340 55168 31248 55196
rect 33060 55196 33088 55236
rect 33134 55224 33140 55276
rect 33192 55264 33198 55276
rect 33229 55267 33287 55273
rect 33229 55264 33241 55267
rect 33192 55236 33241 55264
rect 33192 55224 33198 55236
rect 33229 55233 33241 55236
rect 33275 55233 33287 55267
rect 33229 55227 33287 55233
rect 33594 55224 33600 55276
rect 33652 55264 33658 55276
rect 34716 55273 34744 55304
rect 35434 55292 35440 55344
rect 35492 55332 35498 55344
rect 35492 55304 37412 55332
rect 35492 55292 35498 55304
rect 34701 55267 34759 55273
rect 33652 55236 34652 55264
rect 33652 55224 33658 55236
rect 33689 55199 33747 55205
rect 33689 55196 33701 55199
rect 33060 55168 33701 55196
rect 30340 55156 30346 55168
rect 33689 55165 33701 55168
rect 33735 55165 33747 55199
rect 34624 55196 34652 55236
rect 34701 55233 34713 55267
rect 34747 55233 34759 55267
rect 34701 55227 34759 55233
rect 34977 55267 35035 55273
rect 34977 55233 34989 55267
rect 35023 55264 35035 55267
rect 36170 55264 36176 55276
rect 35023 55236 36176 55264
rect 35023 55233 35035 55236
rect 34977 55227 35035 55233
rect 36170 55224 36176 55236
rect 36228 55224 36234 55276
rect 36814 55224 36820 55276
rect 36872 55264 36878 55276
rect 37274 55264 37280 55276
rect 36872 55236 37280 55264
rect 36872 55224 36878 55236
rect 37274 55224 37280 55236
rect 37332 55224 37338 55276
rect 35529 55199 35587 55205
rect 35529 55196 35541 55199
rect 34624 55168 35541 55196
rect 33689 55159 33747 55165
rect 35529 55165 35541 55168
rect 35575 55165 35587 55199
rect 36262 55196 36268 55208
rect 35529 55159 35587 55165
rect 35636 55168 36268 55196
rect 27249 55131 27307 55137
rect 27249 55097 27261 55131
rect 27295 55128 27307 55131
rect 27614 55128 27620 55140
rect 27295 55100 27620 55128
rect 27295 55097 27307 55100
rect 27249 55091 27307 55097
rect 27614 55088 27620 55100
rect 27672 55088 27678 55140
rect 28258 55128 28264 55140
rect 28219 55100 28264 55128
rect 28258 55088 28264 55100
rect 28316 55088 28322 55140
rect 34793 55131 34851 55137
rect 34793 55097 34805 55131
rect 34839 55097 34851 55131
rect 34793 55091 34851 55097
rect 34885 55131 34943 55137
rect 34885 55097 34897 55131
rect 34931 55128 34943 55131
rect 35636 55128 35664 55168
rect 36262 55156 36268 55168
rect 36320 55156 36326 55208
rect 34931 55100 35664 55128
rect 34931 55097 34943 55100
rect 34885 55091 34943 55097
rect 28445 55063 28503 55069
rect 28445 55029 28457 55063
rect 28491 55060 28503 55063
rect 28718 55060 28724 55072
rect 28491 55032 28724 55060
rect 28491 55029 28503 55032
rect 28445 55023 28503 55029
rect 28718 55020 28724 55032
rect 28776 55020 28782 55072
rect 31846 55020 31852 55072
rect 31904 55060 31910 55072
rect 31941 55063 31999 55069
rect 31941 55060 31953 55063
rect 31904 55032 31953 55060
rect 31904 55020 31910 55032
rect 31941 55029 31953 55032
rect 31987 55029 31999 55063
rect 32306 55060 32312 55072
rect 32267 55032 32312 55060
rect 31941 55023 31999 55029
rect 32306 55020 32312 55032
rect 32364 55020 32370 55072
rect 32766 55060 32772 55072
rect 32727 55032 32772 55060
rect 32766 55020 32772 55032
rect 32824 55020 32830 55072
rect 33137 55063 33195 55069
rect 33137 55029 33149 55063
rect 33183 55060 33195 55063
rect 33410 55060 33416 55072
rect 33183 55032 33416 55060
rect 33183 55029 33195 55032
rect 33137 55023 33195 55029
rect 33410 55020 33416 55032
rect 33468 55020 33474 55072
rect 33870 55020 33876 55072
rect 33928 55060 33934 55072
rect 34808 55060 34836 55091
rect 35986 55088 35992 55140
rect 36044 55128 36050 55140
rect 36173 55131 36231 55137
rect 36173 55128 36185 55131
rect 36044 55100 36185 55128
rect 36044 55088 36050 55100
rect 36173 55097 36185 55100
rect 36219 55097 36231 55131
rect 36173 55091 36231 55097
rect 37277 55131 37335 55137
rect 37277 55097 37289 55131
rect 37323 55128 37335 55131
rect 37384 55128 37412 55304
rect 38746 55292 38752 55344
rect 38804 55332 38810 55344
rect 43070 55332 43076 55344
rect 38804 55304 43076 55332
rect 38804 55292 38810 55304
rect 39040 55273 39068 55304
rect 43070 55292 43076 55304
rect 43128 55292 43134 55344
rect 38197 55267 38255 55273
rect 38197 55233 38209 55267
rect 38243 55264 38255 55267
rect 39025 55267 39083 55273
rect 38243 55236 38976 55264
rect 38243 55233 38255 55236
rect 38197 55227 38255 55233
rect 38381 55199 38439 55205
rect 38381 55165 38393 55199
rect 38427 55196 38439 55199
rect 38746 55196 38752 55208
rect 38427 55168 38752 55196
rect 38427 55165 38439 55168
rect 38381 55159 38439 55165
rect 38746 55156 38752 55168
rect 38804 55156 38810 55208
rect 38948 55196 38976 55236
rect 39025 55233 39037 55267
rect 39071 55233 39083 55267
rect 40218 55264 40224 55276
rect 40131 55236 40224 55264
rect 39025 55227 39083 55233
rect 40218 55224 40224 55236
rect 40276 55224 40282 55276
rect 42061 55267 42119 55273
rect 42061 55233 42073 55267
rect 42107 55264 42119 55267
rect 42518 55264 42524 55276
rect 42107 55236 42524 55264
rect 42107 55233 42119 55236
rect 42061 55227 42119 55233
rect 42518 55224 42524 55236
rect 42576 55224 42582 55276
rect 43165 55267 43223 55273
rect 43165 55233 43177 55267
rect 43211 55264 43223 55267
rect 43898 55264 43904 55276
rect 43211 55236 43904 55264
rect 43211 55233 43223 55236
rect 43165 55227 43223 55233
rect 43898 55224 43904 55236
rect 43956 55224 43962 55276
rect 44008 55273 44036 55372
rect 44358 55360 44364 55372
rect 44416 55360 44422 55412
rect 44726 55400 44732 55412
rect 44687 55372 44732 55400
rect 44726 55360 44732 55372
rect 44784 55360 44790 55412
rect 45554 55400 45560 55412
rect 45515 55372 45560 55400
rect 45554 55360 45560 55372
rect 45612 55360 45618 55412
rect 45646 55360 45652 55412
rect 45704 55400 45710 55412
rect 46109 55403 46167 55409
rect 46109 55400 46121 55403
rect 45704 55372 46121 55400
rect 45704 55360 45710 55372
rect 46109 55369 46121 55372
rect 46155 55369 46167 55403
rect 46109 55363 46167 55369
rect 44266 55292 44272 55344
rect 44324 55332 44330 55344
rect 44324 55304 44956 55332
rect 44324 55292 44330 55304
rect 43993 55267 44051 55273
rect 43993 55233 44005 55267
rect 44039 55233 44051 55267
rect 44174 55264 44180 55276
rect 44135 55236 44180 55264
rect 43993 55227 44051 55233
rect 44174 55224 44180 55236
rect 44232 55224 44238 55276
rect 44928 55273 44956 55304
rect 44913 55267 44971 55273
rect 44913 55233 44925 55267
rect 44959 55233 44971 55267
rect 44913 55227 44971 55233
rect 39117 55199 39175 55205
rect 39117 55196 39129 55199
rect 38948 55168 39129 55196
rect 39117 55165 39129 55168
rect 39163 55165 39175 55199
rect 40236 55196 40264 55224
rect 41969 55199 42027 55205
rect 41969 55196 41981 55199
rect 40236 55168 41981 55196
rect 39117 55159 39175 55165
rect 41969 55165 41981 55168
rect 42015 55196 42027 55199
rect 42610 55196 42616 55208
rect 42015 55168 42616 55196
rect 42015 55165 42027 55168
rect 41969 55159 42027 55165
rect 37323 55100 37412 55128
rect 37323 55097 37335 55100
rect 37277 55091 37335 55097
rect 39022 55088 39028 55140
rect 39080 55128 39086 55140
rect 39132 55128 39160 55159
rect 42610 55156 42616 55168
rect 42668 55196 42674 55208
rect 43257 55199 43315 55205
rect 42668 55168 42932 55196
rect 42668 55156 42674 55168
rect 42797 55131 42855 55137
rect 42797 55128 42809 55131
rect 39080 55100 42809 55128
rect 39080 55088 39086 55100
rect 42797 55097 42809 55100
rect 42843 55097 42855 55131
rect 42904 55128 42932 55168
rect 43257 55165 43269 55199
rect 43303 55196 43315 55199
rect 43809 55199 43867 55205
rect 43809 55196 43821 55199
rect 43303 55168 43821 55196
rect 43303 55165 43315 55168
rect 43257 55159 43315 55165
rect 43809 55165 43821 55168
rect 43855 55165 43867 55199
rect 43809 55159 43867 55165
rect 44082 55156 44088 55208
rect 44140 55196 44146 55208
rect 44269 55199 44327 55205
rect 44269 55196 44281 55199
rect 44140 55168 44281 55196
rect 44140 55156 44146 55168
rect 44269 55165 44281 55168
rect 44315 55165 44327 55199
rect 44269 55159 44327 55165
rect 44100 55128 44128 55156
rect 42904 55100 44128 55128
rect 42797 55091 42855 55097
rect 35710 55060 35716 55072
rect 33928 55032 35716 55060
rect 33928 55020 33934 55032
rect 35710 55020 35716 55032
rect 35768 55020 35774 55072
rect 39393 55063 39451 55069
rect 39393 55029 39405 55063
rect 39439 55060 39451 55063
rect 39666 55060 39672 55072
rect 39439 55032 39672 55060
rect 39439 55029 39451 55032
rect 39393 55023 39451 55029
rect 39666 55020 39672 55032
rect 39724 55020 39730 55072
rect 40497 55063 40555 55069
rect 40497 55029 40509 55063
rect 40543 55060 40555 55063
rect 40586 55060 40592 55072
rect 40543 55032 40592 55060
rect 40543 55029 40555 55032
rect 40497 55023 40555 55029
rect 40586 55020 40592 55032
rect 40644 55020 40650 55072
rect 40681 55063 40739 55069
rect 40681 55029 40693 55063
rect 40727 55060 40739 55063
rect 40770 55060 40776 55072
rect 40727 55032 40776 55060
rect 40727 55029 40739 55032
rect 40681 55023 40739 55029
rect 40770 55020 40776 55032
rect 40828 55020 40834 55072
rect 42242 55060 42248 55072
rect 42203 55032 42248 55060
rect 42242 55020 42248 55032
rect 42300 55020 42306 55072
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 25130 54856 25136 54868
rect 25091 54828 25136 54856
rect 25130 54816 25136 54828
rect 25188 54816 25194 54868
rect 25777 54859 25835 54865
rect 25777 54825 25789 54859
rect 25823 54856 25835 54859
rect 25866 54856 25872 54868
rect 25823 54828 25872 54856
rect 25823 54825 25835 54828
rect 25777 54819 25835 54825
rect 25866 54816 25872 54828
rect 25924 54816 25930 54868
rect 26234 54816 26240 54868
rect 26292 54856 26298 54868
rect 26329 54859 26387 54865
rect 26329 54856 26341 54859
rect 26292 54828 26341 54856
rect 26292 54816 26298 54828
rect 26329 54825 26341 54828
rect 26375 54825 26387 54859
rect 26329 54819 26387 54825
rect 26418 54816 26424 54868
rect 26476 54856 26482 54868
rect 26881 54859 26939 54865
rect 26881 54856 26893 54859
rect 26476 54828 26893 54856
rect 26476 54816 26482 54828
rect 26881 54825 26893 54828
rect 26927 54825 26939 54859
rect 26881 54819 26939 54825
rect 28169 54859 28227 54865
rect 28169 54825 28181 54859
rect 28215 54856 28227 54859
rect 29270 54856 29276 54868
rect 28215 54828 29276 54856
rect 28215 54825 28227 54828
rect 28169 54819 28227 54825
rect 29270 54816 29276 54828
rect 29328 54816 29334 54868
rect 29825 54859 29883 54865
rect 29825 54825 29837 54859
rect 29871 54856 29883 54859
rect 29914 54856 29920 54868
rect 29871 54828 29920 54856
rect 29871 54825 29883 54828
rect 29825 54819 29883 54825
rect 29914 54816 29920 54828
rect 29972 54816 29978 54868
rect 30377 54859 30435 54865
rect 30377 54825 30389 54859
rect 30423 54856 30435 54859
rect 30466 54856 30472 54868
rect 30423 54828 30472 54856
rect 30423 54825 30435 54828
rect 30377 54819 30435 54825
rect 30466 54816 30472 54828
rect 30524 54816 30530 54868
rect 31294 54816 31300 54868
rect 31352 54856 31358 54868
rect 31389 54859 31447 54865
rect 31389 54856 31401 54859
rect 31352 54828 31401 54856
rect 31352 54816 31358 54828
rect 31389 54825 31401 54828
rect 31435 54825 31447 54859
rect 34793 54859 34851 54865
rect 34793 54856 34805 54859
rect 31389 54819 31447 54825
rect 31726 54828 34805 54856
rect 29181 54791 29239 54797
rect 29181 54757 29193 54791
rect 29227 54788 29239 54791
rect 29454 54788 29460 54800
rect 29227 54760 29460 54788
rect 29227 54757 29239 54760
rect 29181 54751 29239 54757
rect 29454 54748 29460 54760
rect 29512 54748 29518 54800
rect 28442 54720 28448 54732
rect 28000 54692 28448 54720
rect 25590 54652 25596 54664
rect 25551 54624 25596 54652
rect 25590 54612 25596 54624
rect 25648 54612 25654 54664
rect 27062 54652 27068 54664
rect 27023 54624 27068 54652
rect 27062 54612 27068 54624
rect 27120 54612 27126 54664
rect 28000 54661 28028 54692
rect 28442 54680 28448 54692
rect 28500 54680 28506 54732
rect 28718 54720 28724 54732
rect 28679 54692 28724 54720
rect 28718 54680 28724 54692
rect 28776 54680 28782 54732
rect 30190 54680 30196 54732
rect 30248 54720 30254 54732
rect 30837 54723 30895 54729
rect 30837 54720 30849 54723
rect 30248 54692 30849 54720
rect 30248 54680 30254 54692
rect 30837 54689 30849 54692
rect 30883 54720 30895 54723
rect 31726 54720 31754 54828
rect 34793 54825 34805 54828
rect 34839 54825 34851 54859
rect 34793 54819 34851 54825
rect 35989 54859 36047 54865
rect 35989 54825 36001 54859
rect 36035 54856 36047 54859
rect 36262 54856 36268 54868
rect 36035 54828 36268 54856
rect 36035 54825 36047 54828
rect 35989 54819 36047 54825
rect 32585 54791 32643 54797
rect 32585 54757 32597 54791
rect 32631 54788 32643 54791
rect 33042 54788 33048 54800
rect 32631 54760 33048 54788
rect 32631 54757 32643 54760
rect 32585 54751 32643 54757
rect 33042 54748 33048 54760
rect 33100 54748 33106 54800
rect 34882 54788 34888 54800
rect 34256 54760 34888 54788
rect 32306 54720 32312 54732
rect 30883 54692 31754 54720
rect 32267 54692 32312 54720
rect 30883 54689 30895 54692
rect 30837 54683 30895 54689
rect 32306 54680 32312 54692
rect 32364 54680 32370 54732
rect 33870 54720 33876 54732
rect 33831 54692 33876 54720
rect 33870 54680 33876 54692
rect 33928 54680 33934 54732
rect 34256 54729 34284 54760
rect 34882 54748 34888 54760
rect 34940 54788 34946 54800
rect 36004 54788 36032 54819
rect 36262 54816 36268 54828
rect 36320 54816 36326 54868
rect 36354 54816 36360 54868
rect 36412 54856 36418 54868
rect 36817 54859 36875 54865
rect 36817 54856 36829 54859
rect 36412 54828 36829 54856
rect 36412 54816 36418 54828
rect 36817 54825 36829 54828
rect 36863 54825 36875 54859
rect 38102 54856 38108 54868
rect 38063 54828 38108 54856
rect 36817 54819 36875 54825
rect 38102 54816 38108 54828
rect 38160 54816 38166 54868
rect 38657 54859 38715 54865
rect 38657 54825 38669 54859
rect 38703 54856 38715 54859
rect 38930 54856 38936 54868
rect 38703 54828 38936 54856
rect 38703 54825 38715 54828
rect 38657 54819 38715 54825
rect 38930 54816 38936 54828
rect 38988 54816 38994 54868
rect 39853 54859 39911 54865
rect 39853 54825 39865 54859
rect 39899 54856 39911 54859
rect 40126 54856 40132 54868
rect 39899 54828 40132 54856
rect 39899 54825 39911 54828
rect 39853 54819 39911 54825
rect 40126 54816 40132 54828
rect 40184 54816 40190 54868
rect 41509 54859 41567 54865
rect 41509 54825 41521 54859
rect 41555 54856 41567 54859
rect 42058 54856 42064 54868
rect 41555 54828 42064 54856
rect 41555 54825 41567 54828
rect 41509 54819 41567 54825
rect 42058 54816 42064 54828
rect 42116 54816 42122 54868
rect 43254 54816 43260 54868
rect 43312 54856 43318 54868
rect 43441 54859 43499 54865
rect 43441 54856 43453 54859
rect 43312 54828 43453 54856
rect 43312 54816 43318 54828
rect 43441 54825 43453 54828
rect 43487 54825 43499 54859
rect 43441 54819 43499 54825
rect 44266 54816 44272 54868
rect 44324 54856 44330 54868
rect 44545 54859 44603 54865
rect 44545 54856 44557 54859
rect 44324 54828 44557 54856
rect 44324 54816 44330 54828
rect 44545 54825 44557 54828
rect 44591 54825 44603 54859
rect 44545 54819 44603 54825
rect 34940 54760 36032 54788
rect 34940 54748 34946 54760
rect 39758 54748 39764 54800
rect 39816 54788 39822 54800
rect 42981 54791 43039 54797
rect 42981 54788 42993 54791
rect 39816 54760 42993 54788
rect 39816 54748 39822 54760
rect 42981 54757 42993 54760
rect 43027 54757 43039 54791
rect 42981 54751 43039 54757
rect 34241 54723 34299 54729
rect 34241 54689 34253 54723
rect 34287 54689 34299 54723
rect 34241 54683 34299 54689
rect 35161 54723 35219 54729
rect 35161 54689 35173 54723
rect 35207 54720 35219 54723
rect 36357 54723 36415 54729
rect 36357 54720 36369 54723
rect 35207 54692 36369 54720
rect 35207 54689 35219 54692
rect 35161 54683 35219 54689
rect 36357 54689 36369 54692
rect 36403 54689 36415 54723
rect 40310 54720 40316 54732
rect 36357 54683 36415 54689
rect 39500 54692 40316 54720
rect 39500 54664 39528 54692
rect 40310 54680 40316 54692
rect 40368 54680 40374 54732
rect 41693 54723 41751 54729
rect 41693 54720 41705 54723
rect 40788 54692 41705 54720
rect 40788 54664 40816 54692
rect 41693 54689 41705 54692
rect 41739 54689 41751 54723
rect 41693 54683 41751 54689
rect 27985 54655 28043 54661
rect 27985 54621 27997 54655
rect 28031 54621 28043 54655
rect 27985 54615 28043 54621
rect 28169 54655 28227 54661
rect 28169 54621 28181 54655
rect 28215 54652 28227 54655
rect 28534 54652 28540 54664
rect 28215 54624 28540 54652
rect 28215 54621 28227 54624
rect 28169 54615 28227 54621
rect 28534 54612 28540 54624
rect 28592 54612 28598 54664
rect 28813 54655 28871 54661
rect 28813 54621 28825 54655
rect 28859 54652 28871 54655
rect 28994 54652 29000 54664
rect 28859 54624 29000 54652
rect 28859 54621 28871 54624
rect 28813 54615 28871 54621
rect 28994 54612 29000 54624
rect 29052 54612 29058 54664
rect 30745 54655 30803 54661
rect 30745 54621 30757 54655
rect 30791 54621 30803 54655
rect 30745 54615 30803 54621
rect 32217 54655 32275 54661
rect 32217 54621 32229 54655
rect 32263 54652 32275 54655
rect 32766 54652 32772 54664
rect 32263 54624 32772 54652
rect 32263 54621 32275 54624
rect 32217 54615 32275 54621
rect 30374 54544 30380 54596
rect 30432 54584 30438 54596
rect 30760 54584 30788 54615
rect 32766 54612 32772 54624
rect 32824 54612 32830 54664
rect 33781 54655 33839 54661
rect 33781 54621 33793 54655
rect 33827 54621 33839 54655
rect 33781 54615 33839 54621
rect 35069 54655 35127 54661
rect 35069 54621 35081 54655
rect 35115 54652 35127 54655
rect 35618 54652 35624 54664
rect 35115 54624 35624 54652
rect 35115 54621 35127 54624
rect 35069 54615 35127 54621
rect 32398 54584 32404 54596
rect 30432 54556 32404 54584
rect 30432 54544 30438 54556
rect 32398 54544 32404 54556
rect 32456 54544 32462 54596
rect 33796 54584 33824 54615
rect 35618 54612 35624 54624
rect 35676 54612 35682 54664
rect 35710 54612 35716 54664
rect 35768 54652 35774 54664
rect 35897 54655 35955 54661
rect 35897 54652 35909 54655
rect 35768 54624 35909 54652
rect 35768 54612 35774 54624
rect 35897 54621 35909 54624
rect 35943 54621 35955 54655
rect 36170 54652 36176 54664
rect 36131 54624 36176 54652
rect 35897 54615 35955 54621
rect 36170 54612 36176 54624
rect 36228 54612 36234 54664
rect 37737 54655 37795 54661
rect 37737 54621 37749 54655
rect 37783 54652 37795 54655
rect 37826 54652 37832 54664
rect 37783 54624 37832 54652
rect 37783 54621 37795 54624
rect 37737 54615 37795 54621
rect 37826 54612 37832 54624
rect 37884 54612 37890 54664
rect 37921 54655 37979 54661
rect 37921 54621 37933 54655
rect 37967 54652 37979 54655
rect 38010 54652 38016 54664
rect 37967 54624 38016 54652
rect 37967 54621 37979 54624
rect 37921 54615 37979 54621
rect 38010 54612 38016 54624
rect 38068 54612 38074 54664
rect 38746 54612 38752 54664
rect 38804 54652 38810 54664
rect 38841 54655 38899 54661
rect 38841 54652 38853 54655
rect 38804 54624 38853 54652
rect 38804 54612 38810 54624
rect 38841 54621 38853 54624
rect 38887 54621 38899 54655
rect 39022 54652 39028 54664
rect 38983 54624 39028 54652
rect 38841 54615 38899 54621
rect 39022 54612 39028 54624
rect 39080 54612 39086 54664
rect 39482 54652 39488 54664
rect 39443 54624 39488 54652
rect 39482 54612 39488 54624
rect 39540 54612 39546 54664
rect 39666 54652 39672 54664
rect 39627 54624 39672 54652
rect 39666 54612 39672 54624
rect 39724 54612 39730 54664
rect 40494 54652 40500 54664
rect 40455 54624 40500 54652
rect 40494 54612 40500 54624
rect 40552 54612 40558 54664
rect 40770 54652 40776 54664
rect 40731 54624 40776 54652
rect 40770 54612 40776 54624
rect 40828 54612 40834 54664
rect 41322 54612 41328 54664
rect 41380 54652 41386 54664
rect 41785 54655 41843 54661
rect 41785 54652 41797 54655
rect 41380 54624 41797 54652
rect 41380 54612 41386 54624
rect 41785 54621 41797 54624
rect 41831 54621 41843 54655
rect 41785 54615 41843 54621
rect 42518 54612 42524 54664
rect 42576 54652 42582 54664
rect 42705 54655 42763 54661
rect 42705 54652 42717 54655
rect 42576 54624 42717 54652
rect 42576 54612 42582 54624
rect 42705 54621 42717 54624
rect 42751 54621 42763 54655
rect 42978 54652 42984 54664
rect 42939 54624 42984 54652
rect 42705 54615 42763 54621
rect 42978 54612 42984 54624
rect 43036 54612 43042 54664
rect 36188 54584 36216 54612
rect 33796 54556 36216 54584
rect 40681 54587 40739 54593
rect 40681 54553 40693 54587
rect 40727 54584 40739 54587
rect 41414 54584 41420 54596
rect 40727 54556 41420 54584
rect 40727 54553 40739 54556
rect 40681 54547 40739 54553
rect 41414 54544 41420 54556
rect 41472 54544 41478 54596
rect 42797 54587 42855 54593
rect 42797 54553 42809 54587
rect 42843 54584 42855 54587
rect 43162 54584 43168 54596
rect 42843 54556 43168 54584
rect 42843 54553 42855 54556
rect 42797 54547 42855 54553
rect 43162 54544 43168 54556
rect 43220 54544 43226 54596
rect 33318 54476 33324 54528
rect 33376 54516 33382 54528
rect 33597 54519 33655 54525
rect 33597 54516 33609 54519
rect 33376 54488 33609 54516
rect 33376 54476 33382 54488
rect 33597 54485 33609 54488
rect 33643 54485 33655 54519
rect 33597 54479 33655 54485
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 26234 54312 26240 54324
rect 26195 54284 26240 54312
rect 26234 54272 26240 54284
rect 26292 54272 26298 54324
rect 29181 54315 29239 54321
rect 29181 54281 29193 54315
rect 29227 54312 29239 54315
rect 29362 54312 29368 54324
rect 29227 54284 29368 54312
rect 29227 54281 29239 54284
rect 29181 54275 29239 54281
rect 29362 54272 29368 54284
rect 29420 54272 29426 54324
rect 30006 54312 30012 54324
rect 29967 54284 30012 54312
rect 30006 54272 30012 54284
rect 30064 54272 30070 54324
rect 30282 54272 30288 54324
rect 30340 54312 30346 54324
rect 31941 54315 31999 54321
rect 31941 54312 31953 54315
rect 30340 54284 31953 54312
rect 30340 54272 30346 54284
rect 31941 54281 31953 54284
rect 31987 54281 31999 54315
rect 31941 54275 31999 54281
rect 32309 54315 32367 54321
rect 32309 54281 32321 54315
rect 32355 54312 32367 54315
rect 32861 54315 32919 54321
rect 32861 54312 32873 54315
rect 32355 54284 32873 54312
rect 32355 54281 32367 54284
rect 32309 54275 32367 54281
rect 32861 54281 32873 54284
rect 32907 54312 32919 54315
rect 33134 54312 33140 54324
rect 32907 54284 33140 54312
rect 32907 54281 32919 54284
rect 32861 54275 32919 54281
rect 33134 54272 33140 54284
rect 33192 54272 33198 54324
rect 33686 54272 33692 54324
rect 33744 54312 33750 54324
rect 33781 54315 33839 54321
rect 33781 54312 33793 54315
rect 33744 54284 33793 54312
rect 33744 54272 33750 54284
rect 33781 54281 33793 54284
rect 33827 54281 33839 54315
rect 33781 54275 33839 54281
rect 36081 54315 36139 54321
rect 36081 54281 36093 54315
rect 36127 54312 36139 54315
rect 36446 54312 36452 54324
rect 36127 54284 36452 54312
rect 36127 54281 36139 54284
rect 36081 54275 36139 54281
rect 36446 54272 36452 54284
rect 36504 54312 36510 54324
rect 36633 54315 36691 54321
rect 36633 54312 36645 54315
rect 36504 54284 36645 54312
rect 36504 54272 36510 54284
rect 36633 54281 36645 54284
rect 36679 54281 36691 54315
rect 36633 54275 36691 54281
rect 39666 54272 39672 54324
rect 39724 54312 39730 54324
rect 40221 54315 40279 54321
rect 40221 54312 40233 54315
rect 39724 54284 40233 54312
rect 39724 54272 39730 54284
rect 40221 54281 40233 54284
rect 40267 54281 40279 54315
rect 41322 54312 41328 54324
rect 41283 54284 41328 54312
rect 40221 54275 40279 54281
rect 41322 54272 41328 54284
rect 41380 54272 41386 54324
rect 41953 54315 42011 54321
rect 41953 54281 41965 54315
rect 41999 54312 42011 54315
rect 42242 54312 42248 54324
rect 41999 54284 42248 54312
rect 41999 54281 42011 54284
rect 41953 54275 42011 54281
rect 42242 54272 42248 54284
rect 42300 54272 42306 54324
rect 42886 54272 42892 54324
rect 42944 54312 42950 54324
rect 43717 54315 43775 54321
rect 43717 54312 43729 54315
rect 42944 54284 43729 54312
rect 42944 54272 42950 54284
rect 43717 54281 43729 54284
rect 43763 54281 43775 54315
rect 43717 54275 43775 54281
rect 29454 54204 29460 54256
rect 29512 54244 29518 54256
rect 29512 54216 30512 54244
rect 29512 54204 29518 54216
rect 26694 54136 26700 54188
rect 26752 54176 26758 54188
rect 26789 54179 26847 54185
rect 26789 54176 26801 54179
rect 26752 54148 26801 54176
rect 26752 54136 26758 54148
rect 26789 54145 26801 54148
rect 26835 54145 26847 54179
rect 26789 54139 26847 54145
rect 28261 54179 28319 54185
rect 28261 54145 28273 54179
rect 28307 54176 28319 54179
rect 28902 54176 28908 54188
rect 28307 54148 28908 54176
rect 28307 54145 28319 54148
rect 28261 54139 28319 54145
rect 28902 54136 28908 54148
rect 28960 54136 28966 54188
rect 29365 54179 29423 54185
rect 29365 54145 29377 54179
rect 29411 54145 29423 54179
rect 29365 54139 29423 54145
rect 29549 54179 29607 54185
rect 29549 54145 29561 54179
rect 29595 54176 29607 54179
rect 30190 54176 30196 54188
rect 29595 54148 30196 54176
rect 29595 54145 29607 54148
rect 29549 54139 29607 54145
rect 29380 54108 29408 54139
rect 30190 54136 30196 54148
rect 30248 54136 30254 54188
rect 30374 54176 30380 54188
rect 30335 54148 30380 54176
rect 30374 54136 30380 54148
rect 30432 54136 30438 54188
rect 30484 54176 30512 54216
rect 30742 54204 30748 54256
rect 30800 54244 30806 54256
rect 30929 54247 30987 54253
rect 30929 54244 30941 54247
rect 30800 54216 30941 54244
rect 30800 54204 30806 54216
rect 30929 54213 30941 54216
rect 30975 54213 30987 54247
rect 33226 54244 33232 54256
rect 33139 54216 33232 54244
rect 30929 54207 30987 54213
rect 33226 54204 33232 54216
rect 33284 54244 33290 54256
rect 34517 54247 34575 54253
rect 34517 54244 34529 54247
rect 33284 54216 34529 54244
rect 33284 54204 33290 54216
rect 34517 54213 34529 54216
rect 34563 54213 34575 54247
rect 36170 54244 36176 54256
rect 34517 54207 34575 54213
rect 34716 54216 36176 54244
rect 30837 54179 30895 54185
rect 30837 54176 30849 54179
rect 30484 54148 30849 54176
rect 30837 54145 30849 54148
rect 30883 54145 30895 54179
rect 31018 54176 31024 54188
rect 30979 54148 31024 54176
rect 30837 54139 30895 54145
rect 31018 54136 31024 54148
rect 31076 54136 31082 54188
rect 32125 54179 32183 54185
rect 32125 54145 32137 54179
rect 32171 54145 32183 54179
rect 32125 54139 32183 54145
rect 30392 54108 30420 54136
rect 29380 54080 30420 54108
rect 32140 54108 32168 54139
rect 32398 54136 32404 54188
rect 32456 54176 32462 54188
rect 32456 54148 32501 54176
rect 32456 54136 32462 54148
rect 32950 54136 32956 54188
rect 33008 54176 33014 54188
rect 33045 54179 33103 54185
rect 33045 54176 33057 54179
rect 33008 54148 33057 54176
rect 33008 54136 33014 54148
rect 33045 54145 33057 54148
rect 33091 54176 33103 54179
rect 33134 54176 33140 54188
rect 33091 54148 33140 54176
rect 33091 54145 33103 54148
rect 33045 54139 33103 54145
rect 33134 54136 33140 54148
rect 33192 54136 33198 54188
rect 33318 54136 33324 54188
rect 33376 54176 33382 54188
rect 33376 54148 33421 54176
rect 33376 54136 33382 54148
rect 33502 54136 33508 54188
rect 33560 54176 33566 54188
rect 33962 54176 33968 54188
rect 33560 54148 33968 54176
rect 33560 54136 33566 54148
rect 33962 54136 33968 54148
rect 34020 54136 34026 54188
rect 34716 54185 34744 54216
rect 36170 54204 36176 54216
rect 36228 54204 36234 54256
rect 40037 54247 40095 54253
rect 40037 54213 40049 54247
rect 40083 54244 40095 54247
rect 40402 54244 40408 54256
rect 40083 54216 40408 54244
rect 40083 54213 40095 54216
rect 40037 54207 40095 54213
rect 40402 54204 40408 54216
rect 40460 54204 40466 54256
rect 41598 54204 41604 54256
rect 41656 54244 41662 54256
rect 42153 54247 42211 54253
rect 42153 54244 42165 54247
rect 41656 54216 42165 54244
rect 41656 54204 41662 54216
rect 42153 54213 42165 54216
rect 42199 54213 42211 54247
rect 42153 54207 42211 54213
rect 34701 54179 34759 54185
rect 34701 54145 34713 54179
rect 34747 54145 34759 54179
rect 34701 54139 34759 54145
rect 34793 54179 34851 54185
rect 34793 54145 34805 54179
rect 34839 54145 34851 54179
rect 34793 54139 34851 54145
rect 33410 54108 33416 54120
rect 32140 54080 33416 54108
rect 33410 54068 33416 54080
rect 33468 54068 33474 54120
rect 34808 54108 34836 54139
rect 34882 54136 34888 54188
rect 34940 54176 34946 54188
rect 34940 54148 34985 54176
rect 34940 54136 34946 54148
rect 35342 54136 35348 54188
rect 35400 54176 35406 54188
rect 35437 54179 35495 54185
rect 35437 54176 35449 54179
rect 35400 54148 35449 54176
rect 35400 54136 35406 54148
rect 35437 54145 35449 54148
rect 35483 54145 35495 54179
rect 37274 54176 37280 54188
rect 37235 54148 37280 54176
rect 35437 54139 35495 54145
rect 37274 54136 37280 54148
rect 37332 54136 37338 54188
rect 37734 54136 37740 54188
rect 37792 54176 37798 54188
rect 37921 54179 37979 54185
rect 37921 54176 37933 54179
rect 37792 54148 37933 54176
rect 37792 54136 37798 54148
rect 37921 54145 37933 54148
rect 37967 54145 37979 54179
rect 37921 54139 37979 54145
rect 38194 54136 38200 54188
rect 38252 54176 38258 54188
rect 38565 54179 38623 54185
rect 38565 54176 38577 54179
rect 38252 54148 38577 54176
rect 38252 54136 38258 54148
rect 38565 54145 38577 54148
rect 38611 54145 38623 54179
rect 38565 54139 38623 54145
rect 39485 54179 39543 54185
rect 39485 54145 39497 54179
rect 39531 54176 39543 54179
rect 39574 54176 39580 54188
rect 39531 54148 39580 54176
rect 39531 54145 39543 54148
rect 39485 54139 39543 54145
rect 39574 54136 39580 54148
rect 39632 54136 39638 54188
rect 40310 54176 40316 54188
rect 40271 54148 40316 54176
rect 40310 54136 40316 54148
rect 40368 54136 40374 54188
rect 40865 54179 40923 54185
rect 40865 54145 40877 54179
rect 40911 54176 40923 54179
rect 41414 54176 41420 54188
rect 40911 54148 41420 54176
rect 40911 54145 40923 54148
rect 40865 54139 40923 54145
rect 41414 54136 41420 54148
rect 41472 54136 41478 54188
rect 42889 54179 42947 54185
rect 42889 54145 42901 54179
rect 42935 54176 42947 54179
rect 43714 54176 43720 54188
rect 42935 54148 43720 54176
rect 42935 54145 42947 54148
rect 42889 54139 42947 54145
rect 43714 54136 43720 54148
rect 43772 54136 43778 54188
rect 35710 54108 35716 54120
rect 34808 54080 35716 54108
rect 35710 54068 35716 54080
rect 35768 54068 35774 54120
rect 28445 54043 28503 54049
rect 28445 54009 28457 54043
rect 28491 54040 28503 54043
rect 31846 54040 31852 54052
rect 28491 54012 31852 54040
rect 28491 54009 28503 54012
rect 28445 54003 28503 54009
rect 31846 54000 31852 54012
rect 31904 54000 31910 54052
rect 40034 54040 40040 54052
rect 39995 54012 40040 54040
rect 40034 54000 40040 54012
rect 40092 54000 40098 54052
rect 27706 53972 27712 53984
rect 27667 53944 27712 53972
rect 27706 53932 27712 53944
rect 27764 53932 27770 53984
rect 40494 53932 40500 53984
rect 40552 53972 40558 53984
rect 40957 53975 41015 53981
rect 40957 53972 40969 53975
rect 40552 53944 40969 53972
rect 40552 53932 40558 53944
rect 40957 53941 40969 53944
rect 41003 53972 41015 53975
rect 41785 53975 41843 53981
rect 41785 53972 41797 53975
rect 41003 53944 41797 53972
rect 41003 53941 41015 53944
rect 40957 53935 41015 53941
rect 41785 53941 41797 53944
rect 41831 53941 41843 53975
rect 41966 53972 41972 53984
rect 41927 53944 41972 53972
rect 41785 53935 41843 53941
rect 41966 53932 41972 53944
rect 42024 53932 42030 53984
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 28074 53768 28080 53780
rect 28035 53740 28080 53768
rect 28074 53728 28080 53740
rect 28132 53728 28138 53780
rect 28629 53771 28687 53777
rect 28629 53737 28641 53771
rect 28675 53768 28687 53771
rect 28902 53768 28908 53780
rect 28675 53740 28908 53768
rect 28675 53737 28687 53740
rect 28629 53731 28687 53737
rect 28902 53728 28908 53740
rect 28960 53728 28966 53780
rect 28994 53728 29000 53780
rect 29052 53768 29058 53780
rect 29641 53771 29699 53777
rect 29641 53768 29653 53771
rect 29052 53740 29653 53768
rect 29052 53728 29058 53740
rect 29641 53737 29653 53740
rect 29687 53737 29699 53771
rect 29641 53731 29699 53737
rect 29730 53728 29736 53780
rect 29788 53768 29794 53780
rect 30377 53771 30435 53777
rect 30377 53768 30389 53771
rect 29788 53740 30389 53768
rect 29788 53728 29794 53740
rect 30377 53737 30389 53740
rect 30423 53737 30435 53771
rect 30377 53731 30435 53737
rect 31018 53728 31024 53780
rect 31076 53768 31082 53780
rect 31113 53771 31171 53777
rect 31113 53768 31125 53771
rect 31076 53740 31125 53768
rect 31076 53728 31082 53740
rect 31113 53737 31125 53740
rect 31159 53737 31171 53771
rect 31938 53768 31944 53780
rect 31899 53740 31944 53768
rect 31113 53731 31171 53737
rect 31938 53728 31944 53740
rect 31996 53728 32002 53780
rect 33226 53728 33232 53780
rect 33284 53768 33290 53780
rect 33321 53771 33379 53777
rect 33321 53768 33333 53771
rect 33284 53740 33333 53768
rect 33284 53728 33290 53740
rect 33321 53737 33333 53740
rect 33367 53737 33379 53771
rect 33962 53768 33968 53780
rect 33923 53740 33968 53768
rect 33321 53731 33379 53737
rect 33962 53728 33968 53740
rect 34020 53728 34026 53780
rect 34790 53728 34796 53780
rect 34848 53768 34854 53780
rect 35069 53771 35127 53777
rect 35069 53768 35081 53771
rect 34848 53740 35081 53768
rect 34848 53728 34854 53740
rect 35069 53737 35081 53740
rect 35115 53737 35127 53771
rect 35069 53731 35127 53737
rect 35989 53771 36047 53777
rect 35989 53737 36001 53771
rect 36035 53768 36047 53771
rect 36078 53768 36084 53780
rect 36035 53740 36084 53768
rect 36035 53737 36047 53740
rect 35989 53731 36047 53737
rect 36078 53728 36084 53740
rect 36136 53768 36142 53780
rect 37001 53771 37059 53777
rect 37001 53768 37013 53771
rect 36136 53740 37013 53768
rect 36136 53728 36142 53740
rect 37001 53737 37013 53740
rect 37047 53737 37059 53771
rect 37001 53731 37059 53737
rect 37458 53728 37464 53780
rect 37516 53768 37522 53780
rect 38657 53771 38715 53777
rect 38657 53768 38669 53771
rect 37516 53740 38669 53768
rect 37516 53728 37522 53740
rect 38657 53737 38669 53740
rect 38703 53737 38715 53771
rect 38657 53731 38715 53737
rect 39393 53771 39451 53777
rect 39393 53737 39405 53771
rect 39439 53768 39451 53771
rect 40402 53768 40408 53780
rect 39439 53740 40408 53768
rect 39439 53737 39451 53740
rect 39393 53731 39451 53737
rect 40402 53728 40408 53740
rect 40460 53768 40466 53780
rect 41417 53771 41475 53777
rect 41417 53768 41429 53771
rect 40460 53740 41429 53768
rect 40460 53728 40466 53740
rect 41417 53737 41429 53740
rect 41463 53768 41475 53771
rect 41969 53771 42027 53777
rect 41969 53768 41981 53771
rect 41463 53740 41981 53768
rect 41463 53737 41475 53740
rect 41417 53731 41475 53737
rect 41969 53737 41981 53740
rect 42015 53737 42027 53771
rect 41969 53731 42027 53737
rect 33137 53703 33195 53709
rect 33137 53669 33149 53703
rect 33183 53700 33195 53703
rect 33410 53700 33416 53712
rect 33183 53672 33416 53700
rect 33183 53669 33195 53672
rect 33137 53663 33195 53669
rect 33410 53660 33416 53672
rect 33468 53660 33474 53712
rect 35894 53660 35900 53712
rect 35952 53700 35958 53712
rect 37553 53703 37611 53709
rect 37553 53700 37565 53703
rect 35952 53672 37565 53700
rect 35952 53660 35958 53672
rect 37553 53669 37565 53672
rect 37599 53669 37611 53703
rect 39850 53700 39856 53712
rect 39811 53672 39856 53700
rect 37553 53663 37611 53669
rect 39850 53660 39856 53672
rect 39908 53660 39914 53712
rect 32582 53632 32588 53644
rect 32495 53604 32588 53632
rect 32582 53592 32588 53604
rect 32640 53632 32646 53644
rect 34609 53635 34667 53641
rect 34609 53632 34621 53635
rect 32640 53604 34621 53632
rect 32640 53592 32646 53604
rect 34609 53601 34621 53604
rect 34655 53632 34667 53635
rect 35986 53632 35992 53644
rect 34655 53604 35992 53632
rect 34655 53601 34667 53604
rect 34609 53595 34667 53601
rect 35986 53592 35992 53604
rect 36044 53632 36050 53644
rect 36446 53632 36452 53644
rect 36044 53604 36452 53632
rect 36044 53592 36050 53604
rect 36446 53592 36452 53604
rect 36504 53592 36510 53644
rect 29178 53524 29184 53576
rect 29236 53564 29242 53576
rect 29365 53567 29423 53573
rect 29365 53564 29377 53567
rect 29236 53536 29377 53564
rect 29236 53524 29242 53536
rect 29365 53533 29377 53536
rect 29411 53533 29423 53567
rect 29365 53527 29423 53533
rect 29641 53567 29699 53573
rect 29641 53533 29653 53567
rect 29687 53564 29699 53567
rect 30006 53564 30012 53576
rect 29687 53536 30012 53564
rect 29687 53533 29699 53536
rect 29641 53527 29699 53533
rect 30006 53524 30012 53536
rect 30064 53524 30070 53576
rect 33134 53524 33140 53576
rect 33192 53564 33198 53576
rect 33192 53536 33548 53564
rect 33192 53524 33198 53536
rect 33318 53505 33324 53508
rect 33305 53499 33324 53505
rect 33305 53465 33317 53499
rect 33305 53459 33324 53465
rect 33318 53456 33324 53459
rect 33376 53456 33382 53508
rect 33520 53505 33548 53536
rect 33505 53499 33563 53505
rect 33505 53465 33517 53499
rect 33551 53465 33563 53499
rect 33505 53459 33563 53465
rect 29362 53388 29368 53440
rect 29420 53428 29426 53440
rect 29457 53431 29515 53437
rect 29457 53428 29469 53431
rect 29420 53400 29469 53428
rect 29420 53388 29426 53400
rect 29457 53397 29469 53400
rect 29503 53397 29515 53431
rect 29457 53391 29515 53397
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 29365 53227 29423 53233
rect 29365 53193 29377 53227
rect 29411 53224 29423 53227
rect 30009 53227 30067 53233
rect 30009 53224 30021 53227
rect 29411 53196 30021 53224
rect 29411 53193 29423 53196
rect 29365 53187 29423 53193
rect 30009 53193 30021 53196
rect 30055 53224 30067 53227
rect 30469 53227 30527 53233
rect 30469 53224 30481 53227
rect 30055 53196 30481 53224
rect 30055 53193 30067 53196
rect 30009 53187 30067 53193
rect 30469 53193 30481 53196
rect 30515 53224 30527 53227
rect 31018 53224 31024 53236
rect 30515 53196 31024 53224
rect 30515 53193 30527 53196
rect 30469 53187 30527 53193
rect 31018 53184 31024 53196
rect 31076 53224 31082 53236
rect 32582 53224 32588 53236
rect 31076 53196 31754 53224
rect 32543 53196 32588 53224
rect 31076 53184 31082 53196
rect 31726 53156 31754 53196
rect 32582 53184 32588 53196
rect 32640 53184 32646 53236
rect 33321 53227 33379 53233
rect 33321 53193 33333 53227
rect 33367 53224 33379 53227
rect 36078 53224 36084 53236
rect 33367 53196 36084 53224
rect 33367 53193 33379 53196
rect 33321 53187 33379 53193
rect 33336 53156 33364 53187
rect 36078 53184 36084 53196
rect 36136 53184 36142 53236
rect 40402 53184 40408 53236
rect 40460 53224 40466 53236
rect 40681 53227 40739 53233
rect 40681 53224 40693 53227
rect 40460 53196 40693 53224
rect 40460 53184 40466 53196
rect 40681 53193 40693 53196
rect 40727 53193 40739 53227
rect 40681 53187 40739 53193
rect 31726 53128 33364 53156
rect 34701 53159 34759 53165
rect 34701 53125 34713 53159
rect 34747 53156 34759 53159
rect 35526 53156 35532 53168
rect 34747 53128 35532 53156
rect 34747 53125 34759 53128
rect 34701 53119 34759 53125
rect 35526 53116 35532 53128
rect 35584 53116 35590 53168
rect 33965 53023 34023 53029
rect 33965 52989 33977 53023
rect 34011 53020 34023 53023
rect 34517 53023 34575 53029
rect 34517 53020 34529 53023
rect 34011 52992 34529 53020
rect 34011 52989 34023 52992
rect 33965 52983 34023 52989
rect 34517 52989 34529 52992
rect 34563 52989 34575 53023
rect 34517 52983 34575 52989
rect 34790 52980 34796 53032
rect 34848 53020 34854 53032
rect 34977 53023 35035 53029
rect 34977 53020 34989 53023
rect 34848 52992 34989 53020
rect 34848 52980 34854 52992
rect 34977 52989 34989 52992
rect 35023 52989 35035 53023
rect 34977 52983 35035 52989
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 35161 52683 35219 52689
rect 35161 52649 35173 52683
rect 35207 52680 35219 52683
rect 35986 52680 35992 52692
rect 35207 52652 35992 52680
rect 35207 52649 35219 52652
rect 35161 52643 35219 52649
rect 35986 52640 35992 52652
rect 36044 52640 36050 52692
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 27706 8032 27712 8084
rect 27764 8072 27770 8084
rect 30653 8075 30711 8081
rect 30653 8072 30665 8075
rect 27764 8044 30665 8072
rect 27764 8032 27770 8044
rect 30653 8041 30665 8044
rect 30699 8072 30711 8075
rect 30834 8072 30840 8084
rect 30699 8044 30840 8072
rect 30699 8041 30711 8044
rect 30653 8035 30711 8041
rect 30834 8032 30840 8044
rect 30892 8072 30898 8084
rect 31573 8075 31631 8081
rect 31573 8072 31585 8075
rect 30892 8044 31585 8072
rect 30892 8032 30898 8044
rect 31573 8041 31585 8044
rect 31619 8041 31631 8075
rect 31573 8035 31631 8041
rect 29549 7871 29607 7877
rect 29549 7837 29561 7871
rect 29595 7868 29607 7871
rect 29638 7868 29644 7880
rect 29595 7840 29644 7868
rect 29595 7837 29607 7840
rect 29549 7831 29607 7837
rect 29638 7828 29644 7840
rect 29696 7828 29702 7880
rect 29457 7735 29515 7741
rect 29457 7701 29469 7735
rect 29503 7732 29515 7735
rect 29546 7732 29552 7744
rect 29503 7704 29552 7732
rect 29503 7701 29515 7704
rect 29457 7695 29515 7701
rect 29546 7692 29552 7704
rect 29604 7692 29610 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 26234 7352 26240 7404
rect 26292 7392 26298 7404
rect 27341 7395 27399 7401
rect 27341 7392 27353 7395
rect 26292 7364 27353 7392
rect 26292 7352 26298 7364
rect 27341 7361 27353 7364
rect 27387 7361 27399 7395
rect 29638 7392 29644 7404
rect 29599 7364 29644 7392
rect 27341 7355 27399 7361
rect 29638 7352 29644 7364
rect 29696 7392 29702 7404
rect 30285 7395 30343 7401
rect 30285 7392 30297 7395
rect 29696 7364 30297 7392
rect 29696 7352 29702 7364
rect 30285 7361 30297 7364
rect 30331 7392 30343 7395
rect 30745 7395 30803 7401
rect 30745 7392 30757 7395
rect 30331 7364 30757 7392
rect 30331 7361 30343 7364
rect 30285 7355 30343 7361
rect 30745 7361 30757 7364
rect 30791 7361 30803 7395
rect 32030 7392 32036 7404
rect 31943 7364 32036 7392
rect 30745 7355 30803 7361
rect 32030 7352 32036 7364
rect 32088 7392 32094 7404
rect 32677 7395 32735 7401
rect 32677 7392 32689 7395
rect 32088 7364 32689 7392
rect 32088 7352 32094 7364
rect 32677 7361 32689 7364
rect 32723 7392 32735 7395
rect 32950 7392 32956 7404
rect 32723 7364 32956 7392
rect 32723 7361 32735 7364
rect 32677 7355 32735 7361
rect 32950 7352 32956 7364
rect 33008 7352 33014 7404
rect 27430 7188 27436 7200
rect 27391 7160 27436 7188
rect 27430 7148 27436 7160
rect 27488 7148 27494 7200
rect 27982 7188 27988 7200
rect 27943 7160 27988 7188
rect 27982 7148 27988 7160
rect 28040 7148 28046 7200
rect 29454 7148 29460 7200
rect 29512 7188 29518 7200
rect 29549 7191 29607 7197
rect 29549 7188 29561 7191
rect 29512 7160 29561 7188
rect 29512 7148 29518 7160
rect 29549 7157 29561 7160
rect 29595 7157 29607 7191
rect 30190 7188 30196 7200
rect 30151 7160 30196 7188
rect 29549 7151 29607 7157
rect 30190 7148 30196 7160
rect 30248 7148 30254 7200
rect 30837 7191 30895 7197
rect 30837 7157 30849 7191
rect 30883 7188 30895 7191
rect 30926 7188 30932 7200
rect 30883 7160 30932 7188
rect 30883 7157 30895 7160
rect 30837 7151 30895 7157
rect 30926 7148 30932 7160
rect 30984 7148 30990 7200
rect 32125 7191 32183 7197
rect 32125 7157 32137 7191
rect 32171 7188 32183 7191
rect 32306 7188 32312 7200
rect 32171 7160 32312 7188
rect 32171 7157 32183 7160
rect 32125 7151 32183 7157
rect 32306 7148 32312 7160
rect 32364 7148 32370 7200
rect 32769 7191 32827 7197
rect 32769 7157 32781 7191
rect 32815 7188 32827 7191
rect 33226 7188 33232 7200
rect 32815 7160 33232 7188
rect 32815 7157 32827 7160
rect 32769 7151 32827 7157
rect 33226 7148 33232 7160
rect 33284 7148 33290 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 31113 6851 31171 6857
rect 31113 6817 31125 6851
rect 31159 6848 31171 6851
rect 32030 6848 32036 6860
rect 31159 6820 32036 6848
rect 31159 6817 31171 6820
rect 31113 6811 31171 6817
rect 32030 6808 32036 6820
rect 32088 6808 32094 6860
rect 25222 6740 25228 6792
rect 25280 6780 25286 6792
rect 25593 6783 25651 6789
rect 25593 6780 25605 6783
rect 25280 6752 25605 6780
rect 25280 6740 25286 6752
rect 25593 6749 25605 6752
rect 25639 6749 25651 6783
rect 26234 6780 26240 6792
rect 26195 6752 26240 6780
rect 25593 6743 25651 6749
rect 26234 6740 26240 6752
rect 26292 6740 26298 6792
rect 26602 6740 26608 6792
rect 26660 6780 26666 6792
rect 26881 6783 26939 6789
rect 26881 6780 26893 6783
rect 26660 6752 26893 6780
rect 26660 6740 26666 6752
rect 26881 6749 26893 6752
rect 26927 6749 26939 6783
rect 27614 6780 27620 6792
rect 27575 6752 27620 6780
rect 26881 6743 26939 6749
rect 27614 6740 27620 6752
rect 27672 6740 27678 6792
rect 28445 6783 28503 6789
rect 28445 6749 28457 6783
rect 28491 6780 28503 6783
rect 28994 6780 29000 6792
rect 28491 6752 29000 6780
rect 28491 6749 28503 6752
rect 28445 6743 28503 6749
rect 28994 6740 29000 6752
rect 29052 6740 29058 6792
rect 29089 6783 29147 6789
rect 29089 6749 29101 6783
rect 29135 6780 29147 6783
rect 29270 6780 29276 6792
rect 29135 6752 29276 6780
rect 29135 6749 29147 6752
rect 29089 6743 29147 6749
rect 29270 6740 29276 6752
rect 29328 6740 29334 6792
rect 29362 6740 29368 6792
rect 29420 6780 29426 6792
rect 29549 6783 29607 6789
rect 29549 6780 29561 6783
rect 29420 6752 29561 6780
rect 29420 6740 29426 6752
rect 29549 6749 29561 6752
rect 29595 6749 29607 6783
rect 30834 6780 30840 6792
rect 30795 6752 30840 6780
rect 29549 6743 29607 6749
rect 30834 6740 30840 6752
rect 30892 6740 30898 6792
rect 31754 6740 31760 6792
rect 31812 6780 31818 6792
rect 32401 6783 32459 6789
rect 31812 6752 31857 6780
rect 31812 6740 31818 6752
rect 32401 6749 32413 6783
rect 32447 6749 32459 6783
rect 33134 6780 33140 6792
rect 33095 6752 33140 6780
rect 32401 6743 32459 6749
rect 29638 6672 29644 6724
rect 29696 6712 29702 6724
rect 32030 6712 32036 6724
rect 29696 6684 32036 6712
rect 29696 6672 29702 6684
rect 32030 6672 32036 6684
rect 32088 6712 32094 6724
rect 32416 6712 32444 6743
rect 33134 6740 33140 6752
rect 33192 6740 33198 6792
rect 33962 6780 33968 6792
rect 33923 6752 33968 6780
rect 33962 6740 33968 6752
rect 34020 6740 34026 6792
rect 32088 6684 32444 6712
rect 32088 6672 32094 6684
rect 25130 6644 25136 6656
rect 25091 6616 25136 6644
rect 25130 6604 25136 6616
rect 25188 6604 25194 6656
rect 26329 6647 26387 6653
rect 26329 6613 26341 6647
rect 26375 6644 26387 6647
rect 26786 6644 26792 6656
rect 26375 6616 26792 6644
rect 26375 6613 26387 6616
rect 26329 6607 26387 6613
rect 26786 6604 26792 6616
rect 26844 6604 26850 6656
rect 32493 6647 32551 6653
rect 32493 6613 32505 6647
rect 32539 6644 32551 6647
rect 33410 6644 33416 6656
rect 32539 6616 33416 6644
rect 32539 6613 32551 6616
rect 32493 6607 32551 6613
rect 33410 6604 33416 6616
rect 33468 6604 33474 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 25041 6443 25099 6449
rect 25041 6409 25053 6443
rect 25087 6440 25099 6443
rect 25130 6440 25136 6452
rect 25087 6412 25136 6440
rect 25087 6409 25099 6412
rect 25041 6403 25099 6409
rect 25130 6400 25136 6412
rect 25188 6440 25194 6452
rect 27706 6440 27712 6452
rect 25188 6412 27712 6440
rect 25188 6400 25194 6412
rect 25700 6316 25728 6412
rect 27706 6400 27712 6412
rect 27764 6400 27770 6452
rect 26786 6372 26792 6384
rect 26747 6344 26792 6372
rect 26786 6332 26792 6344
rect 26844 6332 26850 6384
rect 29454 6372 29460 6384
rect 29415 6344 29460 6372
rect 29454 6332 29460 6344
rect 29512 6332 29518 6384
rect 32030 6372 32036 6384
rect 31991 6344 32036 6372
rect 32030 6332 32036 6344
rect 32088 6332 32094 6384
rect 25682 6304 25688 6316
rect 25595 6276 25688 6304
rect 25682 6264 25688 6276
rect 25740 6264 25746 6316
rect 29270 6304 29276 6316
rect 29231 6276 29276 6304
rect 29270 6264 29276 6276
rect 29328 6264 29334 6316
rect 30834 6264 30840 6316
rect 30892 6304 30898 6316
rect 31757 6307 31815 6313
rect 31757 6304 31769 6307
rect 30892 6276 31769 6304
rect 30892 6264 30898 6276
rect 31757 6273 31769 6276
rect 31803 6273 31815 6307
rect 31757 6267 31815 6273
rect 32950 6264 32956 6316
rect 33008 6304 33014 6316
rect 34517 6307 34575 6313
rect 34517 6304 34529 6307
rect 33008 6276 34529 6304
rect 33008 6264 33014 6276
rect 34517 6273 34529 6276
rect 34563 6273 34575 6307
rect 34517 6267 34575 6273
rect 24854 6196 24860 6248
rect 24912 6236 24918 6248
rect 26605 6239 26663 6245
rect 26605 6236 26617 6239
rect 24912 6208 26617 6236
rect 24912 6196 24918 6208
rect 26605 6205 26617 6208
rect 26651 6205 26663 6239
rect 27522 6236 27528 6248
rect 27483 6208 27528 6236
rect 26605 6199 26663 6205
rect 27522 6196 27528 6208
rect 27580 6196 27586 6248
rect 30006 6236 30012 6248
rect 29967 6208 30012 6236
rect 30006 6196 30012 6208
rect 30064 6196 30070 6248
rect 32861 6171 32919 6177
rect 32861 6137 32873 6171
rect 32907 6168 32919 6171
rect 33594 6168 33600 6180
rect 32907 6140 33600 6168
rect 32907 6137 32919 6140
rect 32861 6131 32919 6137
rect 33594 6128 33600 6140
rect 33652 6128 33658 6180
rect 25406 6060 25412 6112
rect 25464 6100 25470 6112
rect 25593 6103 25651 6109
rect 25593 6100 25605 6103
rect 25464 6072 25605 6100
rect 25464 6060 25470 6072
rect 25593 6069 25605 6072
rect 25639 6069 25651 6103
rect 25593 6063 25651 6069
rect 32122 6060 32128 6112
rect 32180 6100 32186 6112
rect 33321 6103 33379 6109
rect 33321 6100 33333 6103
rect 32180 6072 33333 6100
rect 32180 6060 32186 6072
rect 33321 6069 33333 6072
rect 33367 6069 33379 6103
rect 33321 6063 33379 6069
rect 34609 6103 34667 6109
rect 34609 6069 34621 6103
rect 34655 6100 34667 6103
rect 34790 6100 34796 6112
rect 34655 6072 34796 6100
rect 34655 6069 34667 6072
rect 34609 6063 34667 6069
rect 34790 6060 34796 6072
rect 34848 6060 34854 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 31754 5828 31760 5840
rect 30760 5800 31760 5828
rect 26694 5760 26700 5772
rect 26655 5732 26700 5760
rect 26694 5720 26700 5732
rect 26752 5720 26758 5772
rect 28626 5760 28632 5772
rect 28587 5732 28632 5760
rect 28626 5720 28632 5732
rect 28684 5720 28690 5772
rect 30760 5769 30788 5800
rect 31754 5788 31760 5800
rect 31812 5788 31818 5840
rect 33962 5788 33968 5840
rect 34020 5828 34026 5840
rect 34020 5800 35020 5828
rect 34020 5788 34026 5800
rect 30745 5763 30803 5769
rect 30745 5729 30757 5763
rect 30791 5729 30803 5763
rect 30926 5760 30932 5772
rect 30887 5732 30932 5760
rect 30745 5723 30803 5729
rect 30926 5720 30932 5732
rect 30984 5720 30990 5772
rect 31662 5760 31668 5772
rect 31623 5732 31668 5760
rect 31662 5720 31668 5732
rect 31720 5720 31726 5772
rect 33318 5760 33324 5772
rect 33279 5732 33324 5760
rect 33318 5720 33324 5732
rect 33376 5720 33382 5772
rect 34790 5760 34796 5772
rect 34751 5732 34796 5760
rect 34790 5720 34796 5732
rect 34848 5720 34854 5772
rect 34992 5769 35020 5800
rect 34977 5763 35035 5769
rect 34977 5729 34989 5763
rect 35023 5729 35035 5763
rect 34977 5723 35035 5729
rect 23382 5652 23388 5704
rect 23440 5692 23446 5704
rect 23477 5695 23535 5701
rect 23477 5692 23489 5695
rect 23440 5664 23489 5692
rect 23440 5652 23446 5664
rect 23477 5661 23489 5664
rect 23523 5661 23535 5695
rect 24302 5692 24308 5704
rect 24263 5664 24308 5692
rect 23477 5655 23535 5661
rect 24302 5652 24308 5664
rect 24360 5652 24366 5704
rect 24946 5652 24952 5704
rect 25004 5692 25010 5704
rect 25225 5695 25283 5701
rect 25225 5692 25237 5695
rect 25004 5664 25237 5692
rect 25004 5652 25010 5664
rect 25225 5661 25237 5664
rect 25271 5661 25283 5695
rect 27890 5692 27896 5704
rect 27851 5664 27896 5692
rect 25225 5655 25283 5661
rect 27890 5652 27896 5664
rect 27948 5652 27954 5704
rect 25409 5627 25467 5633
rect 25409 5593 25421 5627
rect 25455 5624 25467 5627
rect 25498 5624 25504 5636
rect 25455 5596 25504 5624
rect 25455 5593 25467 5596
rect 25409 5587 25467 5593
rect 25498 5584 25504 5596
rect 25556 5584 25562 5636
rect 28074 5624 28080 5636
rect 28035 5596 28080 5624
rect 28074 5584 28080 5596
rect 28132 5584 28138 5636
rect 24026 5516 24032 5568
rect 24084 5556 24090 5568
rect 24213 5559 24271 5565
rect 24213 5556 24225 5559
rect 24084 5528 24225 5556
rect 24084 5516 24090 5528
rect 24213 5525 24225 5528
rect 24259 5525 24271 5559
rect 24213 5519 24271 5525
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 25409 5287 25467 5293
rect 25409 5253 25421 5287
rect 25455 5284 25467 5287
rect 26142 5284 26148 5296
rect 25455 5256 26148 5284
rect 25455 5253 25467 5256
rect 25409 5247 25467 5253
rect 24302 5176 24308 5228
rect 24360 5216 24366 5228
rect 24581 5219 24639 5225
rect 24581 5216 24593 5219
rect 24360 5188 24593 5216
rect 24360 5176 24366 5188
rect 24581 5185 24593 5188
rect 24627 5216 24639 5219
rect 25424 5216 25452 5247
rect 26142 5244 26148 5256
rect 26200 5244 26206 5296
rect 26789 5287 26847 5293
rect 26789 5253 26801 5287
rect 26835 5284 26847 5287
rect 27430 5284 27436 5296
rect 26835 5256 27436 5284
rect 26835 5253 26847 5256
rect 26789 5247 26847 5253
rect 27430 5244 27436 5256
rect 27488 5244 27494 5296
rect 29549 5287 29607 5293
rect 29549 5253 29561 5287
rect 29595 5284 29607 5287
rect 30190 5284 30196 5296
rect 29595 5256 30196 5284
rect 29595 5253 29607 5256
rect 29549 5247 29607 5253
rect 30190 5244 30196 5256
rect 30248 5244 30254 5296
rect 33410 5284 33416 5296
rect 33371 5256 33416 5284
rect 33410 5244 33416 5256
rect 33468 5244 33474 5296
rect 36173 5287 36231 5293
rect 36173 5253 36185 5287
rect 36219 5284 36231 5287
rect 37918 5284 37924 5296
rect 36219 5256 37924 5284
rect 36219 5253 36231 5256
rect 36173 5247 36231 5253
rect 37918 5244 37924 5256
rect 37976 5244 37982 5296
rect 25682 5216 25688 5228
rect 24627 5188 25452 5216
rect 25643 5188 25688 5216
rect 24627 5185 24639 5188
rect 24581 5179 24639 5185
rect 25682 5176 25688 5188
rect 25740 5176 25746 5228
rect 26602 5216 26608 5228
rect 26563 5188 26608 5216
rect 26602 5176 26608 5188
rect 26660 5176 26666 5228
rect 29362 5216 29368 5228
rect 29323 5188 29368 5216
rect 29362 5176 29368 5188
rect 29420 5176 29426 5228
rect 33594 5176 33600 5228
rect 33652 5216 33658 5228
rect 33652 5188 33697 5216
rect 33652 5176 33658 5188
rect 24121 5151 24179 5157
rect 24121 5117 24133 5151
rect 24167 5148 24179 5151
rect 24854 5148 24860 5160
rect 24167 5120 24860 5148
rect 24167 5117 24179 5120
rect 24121 5111 24179 5117
rect 24854 5108 24860 5120
rect 24912 5108 24918 5160
rect 27706 5148 27712 5160
rect 27667 5120 27712 5148
rect 27706 5108 27712 5120
rect 27764 5108 27770 5160
rect 30374 5148 30380 5160
rect 30335 5120 30380 5148
rect 30374 5108 30380 5120
rect 30432 5108 30438 5160
rect 31754 5108 31760 5160
rect 31812 5148 31818 5160
rect 34514 5148 34520 5160
rect 31812 5120 31857 5148
rect 34475 5120 34520 5148
rect 31812 5108 31818 5120
rect 34514 5108 34520 5120
rect 34572 5108 34578 5160
rect 36357 5151 36415 5157
rect 36357 5117 36369 5151
rect 36403 5148 36415 5151
rect 37182 5148 37188 5160
rect 36403 5120 37188 5148
rect 36403 5117 36415 5120
rect 36357 5111 36415 5117
rect 37182 5108 37188 5120
rect 37240 5108 37246 5160
rect 22554 4972 22560 5024
rect 22612 5012 22618 5024
rect 22649 5015 22707 5021
rect 22649 5012 22661 5015
rect 22612 4984 22661 5012
rect 22612 4972 22618 4984
rect 22649 4981 22661 4984
rect 22695 4981 22707 5015
rect 22649 4975 22707 4981
rect 24673 5015 24731 5021
rect 24673 4981 24685 5015
rect 24719 5012 24731 5015
rect 27798 5012 27804 5024
rect 24719 4984 27804 5012
rect 24719 4981 24731 4984
rect 24673 4975 24731 4981
rect 27798 4972 27804 4984
rect 27856 4972 27862 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 37182 4808 37188 4820
rect 37143 4780 37188 4808
rect 37182 4768 37188 4780
rect 37240 4768 37246 4820
rect 22373 4743 22431 4749
rect 22373 4709 22385 4743
rect 22419 4740 22431 4743
rect 23934 4740 23940 4752
rect 22419 4712 23940 4740
rect 22419 4709 22431 4712
rect 22373 4703 22431 4709
rect 23934 4700 23940 4712
rect 23992 4700 23998 4752
rect 33226 4700 33232 4752
rect 33284 4740 33290 4752
rect 33284 4712 33364 4740
rect 33284 4700 33290 4712
rect 23661 4675 23719 4681
rect 23661 4641 23673 4675
rect 23707 4672 23719 4675
rect 25038 4672 25044 4684
rect 23707 4644 25044 4672
rect 23707 4641 23719 4644
rect 23661 4635 23719 4641
rect 25038 4632 25044 4644
rect 25096 4632 25102 4684
rect 25222 4672 25228 4684
rect 25183 4644 25228 4672
rect 25222 4632 25228 4644
rect 25280 4632 25286 4684
rect 25406 4672 25412 4684
rect 25367 4644 25412 4672
rect 25406 4632 25412 4644
rect 25464 4632 25470 4684
rect 26234 4672 26240 4684
rect 26195 4644 26240 4672
rect 26234 4632 26240 4644
rect 26292 4632 26298 4684
rect 27614 4672 27620 4684
rect 27575 4644 27620 4672
rect 27614 4632 27620 4644
rect 27672 4632 27678 4684
rect 27798 4672 27804 4684
rect 27759 4644 27804 4672
rect 27798 4632 27804 4644
rect 27856 4632 27862 4684
rect 28166 4672 28172 4684
rect 28127 4644 28172 4672
rect 28166 4632 28172 4644
rect 28224 4632 28230 4684
rect 30742 4632 30748 4684
rect 30800 4672 30806 4684
rect 30837 4675 30895 4681
rect 30837 4672 30849 4675
rect 30800 4644 30849 4672
rect 30800 4632 30806 4644
rect 30837 4641 30849 4644
rect 30883 4641 30895 4675
rect 33134 4672 33140 4684
rect 33095 4644 33140 4672
rect 30837 4635 30895 4641
rect 33134 4632 33140 4644
rect 33192 4632 33198 4684
rect 33336 4681 33364 4712
rect 33321 4675 33379 4681
rect 33321 4641 33333 4675
rect 33367 4641 33379 4675
rect 33594 4672 33600 4684
rect 33555 4644 33600 4672
rect 33321 4635 33379 4641
rect 33594 4632 33600 4644
rect 33652 4632 33658 4684
rect 20714 4604 20720 4616
rect 20675 4576 20720 4604
rect 20714 4564 20720 4576
rect 20772 4564 20778 4616
rect 21545 4607 21603 4613
rect 21545 4573 21557 4607
rect 21591 4604 21603 4607
rect 22002 4604 22008 4616
rect 21591 4576 22008 4604
rect 21591 4573 21603 4576
rect 21545 4567 21603 4573
rect 22002 4564 22008 4576
rect 22060 4564 22066 4616
rect 23017 4607 23075 4613
rect 23017 4573 23029 4607
rect 23063 4604 23075 4607
rect 23474 4604 23480 4616
rect 23063 4576 23480 4604
rect 23063 4573 23075 4576
rect 23017 4567 23075 4573
rect 23474 4564 23480 4576
rect 23532 4604 23538 4616
rect 24121 4607 24179 4613
rect 24121 4604 24133 4607
rect 23532 4576 24133 4604
rect 23532 4564 23538 4576
rect 24121 4573 24133 4576
rect 24167 4604 24179 4607
rect 24302 4604 24308 4616
rect 24167 4576 24308 4604
rect 24167 4573 24179 4576
rect 24121 4567 24179 4573
rect 24302 4564 24308 4576
rect 24360 4564 24366 4616
rect 30374 4604 30380 4616
rect 30335 4576 30380 4604
rect 30374 4564 30380 4576
rect 30432 4564 30438 4616
rect 36081 4607 36139 4613
rect 36081 4573 36093 4607
rect 36127 4604 36139 4607
rect 36354 4604 36360 4616
rect 36127 4576 36360 4604
rect 36127 4573 36139 4576
rect 36081 4567 36139 4573
rect 36354 4564 36360 4576
rect 36412 4564 36418 4616
rect 36722 4604 36728 4616
rect 36683 4576 36728 4604
rect 36722 4564 36728 4576
rect 36780 4564 36786 4616
rect 37826 4604 37832 4616
rect 37787 4576 37832 4604
rect 37826 4564 37832 4576
rect 37884 4564 37890 4616
rect 30561 4539 30619 4545
rect 30561 4505 30573 4539
rect 30607 4536 30619 4539
rect 30650 4536 30656 4548
rect 30607 4508 30656 4536
rect 30607 4505 30619 4508
rect 30561 4499 30619 4505
rect 30650 4496 30656 4508
rect 30708 4496 30714 4548
rect 22646 4428 22652 4480
rect 22704 4468 22710 4480
rect 22925 4471 22983 4477
rect 22925 4468 22937 4471
rect 22704 4440 22937 4468
rect 22704 4428 22710 4440
rect 22925 4437 22937 4440
rect 22971 4437 22983 4471
rect 22925 4431 22983 4437
rect 24213 4471 24271 4477
rect 24213 4437 24225 4471
rect 24259 4468 24271 4471
rect 26142 4468 26148 4480
rect 24259 4440 26148 4468
rect 24259 4437 24271 4440
rect 24213 4431 24271 4437
rect 26142 4428 26148 4440
rect 26200 4428 26206 4480
rect 36170 4428 36176 4480
rect 36228 4468 36234 4480
rect 36633 4471 36691 4477
rect 36633 4468 36645 4471
rect 36228 4440 36645 4468
rect 36228 4428 36234 4440
rect 36633 4437 36645 4440
rect 36679 4437 36691 4471
rect 36633 4431 36691 4437
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 36170 4196 36176 4208
rect 36131 4168 36176 4196
rect 36170 4156 36176 4168
rect 36228 4156 36234 4208
rect 22741 4131 22799 4137
rect 22741 4097 22753 4131
rect 22787 4128 22799 4131
rect 23474 4128 23480 4140
rect 22787 4100 23480 4128
rect 22787 4097 22799 4100
rect 22741 4091 22799 4097
rect 23474 4088 23480 4100
rect 23532 4088 23538 4140
rect 25314 4088 25320 4140
rect 25372 4128 25378 4140
rect 26605 4131 26663 4137
rect 26605 4128 26617 4131
rect 25372 4100 26617 4128
rect 25372 4088 25378 4100
rect 26605 4097 26617 4100
rect 26651 4097 26663 4131
rect 26605 4091 26663 4097
rect 28994 4088 29000 4140
rect 29052 4128 29058 4140
rect 29181 4131 29239 4137
rect 29181 4128 29193 4131
rect 29052 4100 29193 4128
rect 29052 4088 29058 4100
rect 29181 4097 29193 4100
rect 29227 4097 29239 4131
rect 32122 4128 32128 4140
rect 32083 4100 32128 4128
rect 29181 4091 29239 4097
rect 32122 4088 32128 4100
rect 32180 4088 32186 4140
rect 36354 4088 36360 4140
rect 36412 4128 36418 4140
rect 36412 4100 36457 4128
rect 36412 4088 36418 4100
rect 20993 4063 21051 4069
rect 20993 4029 21005 4063
rect 21039 4060 21051 4063
rect 22278 4060 22284 4072
rect 21039 4032 22284 4060
rect 21039 4029 21051 4032
rect 20993 4023 21051 4029
rect 22278 4020 22284 4032
rect 22336 4020 22342 4072
rect 23842 4060 23848 4072
rect 23803 4032 23848 4060
rect 23842 4020 23848 4032
rect 23900 4020 23906 4072
rect 24029 4063 24087 4069
rect 24029 4029 24041 4063
rect 24075 4029 24087 4063
rect 24029 4023 24087 4029
rect 25685 4063 25743 4069
rect 25685 4029 25697 4063
rect 25731 4029 25743 4063
rect 25685 4023 25743 4029
rect 26789 4063 26847 4069
rect 26789 4029 26801 4063
rect 26835 4029 26847 4063
rect 26789 4023 26847 4029
rect 28445 4063 28503 4069
rect 28445 4029 28457 4063
rect 28491 4060 28503 4063
rect 29365 4063 29423 4069
rect 28491 4032 29224 4060
rect 28491 4029 28503 4032
rect 28445 4023 28503 4029
rect 21637 3995 21695 4001
rect 21637 3961 21649 3995
rect 21683 3992 21695 3995
rect 22094 3992 22100 4004
rect 21683 3964 22100 3992
rect 21683 3961 21695 3964
rect 21637 3955 21695 3961
rect 22094 3952 22100 3964
rect 22152 3952 22158 4004
rect 22186 3952 22192 4004
rect 22244 3992 22250 4004
rect 24044 3992 24072 4023
rect 22244 3964 24072 3992
rect 22244 3952 22250 3964
rect 17126 3884 17132 3936
rect 17184 3924 17190 3936
rect 17221 3927 17279 3933
rect 17221 3924 17233 3927
rect 17184 3896 17233 3924
rect 17184 3884 17190 3896
rect 17221 3893 17233 3896
rect 17267 3893 17279 3927
rect 17221 3887 17279 3893
rect 18414 3884 18420 3936
rect 18472 3924 18478 3936
rect 18509 3927 18567 3933
rect 18509 3924 18521 3927
rect 18472 3896 18521 3924
rect 18472 3884 18478 3896
rect 18509 3893 18521 3896
rect 18555 3893 18567 3927
rect 18509 3887 18567 3893
rect 19521 3927 19579 3933
rect 19521 3893 19533 3927
rect 19567 3924 19579 3927
rect 20070 3924 20076 3936
rect 19567 3896 20076 3924
rect 19567 3893 19579 3896
rect 19521 3887 19579 3893
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20165 3927 20223 3933
rect 20165 3893 20177 3927
rect 20211 3924 20223 3927
rect 20346 3924 20352 3936
rect 20211 3896 20352 3924
rect 20211 3893 20223 3896
rect 20165 3887 20223 3893
rect 20346 3884 20352 3896
rect 20404 3884 20410 3936
rect 22281 3927 22339 3933
rect 22281 3893 22293 3927
rect 22327 3924 22339 3927
rect 22462 3924 22468 3936
rect 22327 3896 22468 3924
rect 22327 3893 22339 3896
rect 22281 3887 22339 3893
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 22833 3927 22891 3933
rect 22833 3893 22845 3927
rect 22879 3924 22891 3927
rect 25130 3924 25136 3936
rect 22879 3896 25136 3924
rect 22879 3893 22891 3896
rect 22833 3887 22891 3893
rect 25130 3884 25136 3896
rect 25188 3884 25194 3936
rect 25700 3924 25728 4023
rect 26510 3952 26516 4004
rect 26568 3992 26574 4004
rect 26804 3992 26832 4023
rect 29196 4004 29224 4032
rect 29365 4029 29377 4063
rect 29411 4060 29423 4063
rect 29546 4060 29552 4072
rect 29411 4032 29552 4060
rect 29411 4029 29423 4032
rect 29365 4023 29423 4029
rect 29546 4020 29552 4032
rect 29604 4020 29610 4072
rect 29730 4060 29736 4072
rect 29691 4032 29736 4060
rect 29730 4020 29736 4032
rect 29788 4020 29794 4072
rect 32306 4060 32312 4072
rect 32267 4032 32312 4060
rect 32306 4020 32312 4032
rect 32364 4020 32370 4072
rect 32766 4060 32772 4072
rect 32727 4032 32772 4060
rect 32766 4020 32772 4032
rect 32824 4020 32830 4072
rect 34054 4020 34060 4072
rect 34112 4060 34118 4072
rect 34517 4063 34575 4069
rect 34517 4060 34529 4063
rect 34112 4032 34529 4060
rect 34112 4020 34118 4032
rect 34517 4029 34529 4032
rect 34563 4029 34575 4063
rect 34517 4023 34575 4029
rect 35802 4020 35808 4072
rect 35860 4060 35866 4072
rect 37921 4063 37979 4069
rect 37921 4060 37933 4063
rect 35860 4032 37933 4060
rect 35860 4020 35866 4032
rect 37921 4029 37933 4032
rect 37967 4029 37979 4063
rect 37921 4023 37979 4029
rect 39114 4020 39120 4072
rect 39172 4060 39178 4072
rect 40037 4063 40095 4069
rect 40037 4060 40049 4063
rect 39172 4032 40049 4060
rect 39172 4020 39178 4032
rect 40037 4029 40049 4032
rect 40083 4029 40095 4063
rect 40037 4023 40095 4029
rect 26568 3964 26832 3992
rect 26568 3952 26574 3964
rect 29178 3952 29184 4004
rect 29236 3952 29242 4004
rect 37550 3952 37556 4004
rect 37608 3992 37614 4004
rect 38565 3995 38623 4001
rect 38565 3992 38577 3995
rect 37608 3964 38577 3992
rect 37608 3952 37614 3964
rect 38565 3961 38577 3964
rect 38611 3961 38623 3995
rect 38565 3955 38623 3961
rect 39942 3952 39948 4004
rect 40000 3992 40006 4004
rect 40681 3995 40739 4001
rect 40681 3992 40693 3995
rect 40000 3964 40693 3992
rect 40000 3952 40006 3964
rect 40681 3961 40693 3964
rect 40727 3961 40739 3995
rect 40681 3955 40739 3961
rect 26970 3924 26976 3936
rect 25700 3896 26976 3924
rect 26970 3884 26976 3896
rect 27028 3884 27034 3936
rect 37274 3924 37280 3936
rect 37235 3896 37280 3924
rect 37274 3884 37280 3896
rect 37332 3884 37338 3936
rect 38286 3884 38292 3936
rect 38344 3924 38350 3936
rect 39209 3927 39267 3933
rect 39209 3924 39221 3927
rect 38344 3896 39221 3924
rect 38344 3884 38350 3896
rect 39209 3893 39221 3896
rect 39255 3893 39267 3927
rect 39209 3887 39267 3893
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 22094 3680 22100 3732
rect 22152 3720 22158 3732
rect 24946 3720 24952 3732
rect 22152 3692 24952 3720
rect 22152 3680 22158 3692
rect 24946 3680 24952 3692
rect 25004 3680 25010 3732
rect 25130 3680 25136 3732
rect 25188 3720 25194 3732
rect 28074 3720 28080 3732
rect 25188 3692 28080 3720
rect 25188 3680 25194 3692
rect 28074 3680 28080 3692
rect 28132 3680 28138 3732
rect 36906 3680 36912 3732
rect 36964 3720 36970 3732
rect 37826 3720 37832 3732
rect 36964 3692 37832 3720
rect 36964 3680 36970 3692
rect 37826 3680 37832 3692
rect 37884 3680 37890 3732
rect 20257 3655 20315 3661
rect 20257 3621 20269 3655
rect 20303 3652 20315 3655
rect 21726 3652 21732 3664
rect 20303 3624 21732 3652
rect 20303 3621 20315 3624
rect 20257 3615 20315 3621
rect 21726 3612 21732 3624
rect 21784 3612 21790 3664
rect 26142 3612 26148 3664
rect 26200 3652 26206 3664
rect 26200 3624 28212 3652
rect 26200 3612 26206 3624
rect 19613 3587 19671 3593
rect 19613 3553 19625 3587
rect 19659 3584 19671 3587
rect 21174 3584 21180 3596
rect 19659 3556 21180 3584
rect 19659 3553 19671 3556
rect 19613 3547 19671 3553
rect 21174 3544 21180 3556
rect 21232 3544 21238 3596
rect 22462 3584 22468 3596
rect 22423 3556 22468 3584
rect 22462 3544 22468 3556
rect 22520 3544 22526 3596
rect 22646 3584 22652 3596
rect 22607 3556 22652 3584
rect 22646 3544 22652 3556
rect 22704 3544 22710 3596
rect 25038 3544 25044 3596
rect 25096 3584 25102 3596
rect 25225 3587 25283 3593
rect 25225 3584 25237 3587
rect 25096 3556 25237 3584
rect 25096 3544 25102 3556
rect 25225 3553 25237 3556
rect 25271 3553 25283 3587
rect 27982 3584 27988 3596
rect 27943 3556 27988 3584
rect 25225 3547 25283 3553
rect 27982 3544 27988 3556
rect 28040 3544 28046 3596
rect 28184 3593 28212 3624
rect 36170 3612 36176 3664
rect 36228 3652 36234 3664
rect 38657 3655 38715 3661
rect 38657 3652 38669 3655
rect 36228 3624 38669 3652
rect 36228 3612 36234 3624
rect 38657 3621 38669 3624
rect 38703 3621 38715 3655
rect 38657 3615 38715 3621
rect 40494 3612 40500 3664
rect 40552 3652 40558 3664
rect 41417 3655 41475 3661
rect 41417 3652 41429 3655
rect 40552 3624 41429 3652
rect 40552 3612 40558 3624
rect 41417 3621 41429 3624
rect 41463 3621 41475 3655
rect 41417 3615 41475 3621
rect 42702 3612 42708 3664
rect 42760 3652 42766 3664
rect 43349 3655 43407 3661
rect 43349 3652 43361 3655
rect 42760 3624 43361 3652
rect 42760 3612 42766 3624
rect 43349 3621 43361 3624
rect 43395 3621 43407 3655
rect 43349 3615 43407 3621
rect 28169 3587 28227 3593
rect 28169 3553 28181 3587
rect 28215 3553 28227 3587
rect 28169 3547 28227 3553
rect 28350 3544 28356 3596
rect 28408 3584 28414 3596
rect 28445 3587 28503 3593
rect 28445 3584 28457 3587
rect 28408 3556 28457 3584
rect 28408 3544 28414 3556
rect 28445 3553 28457 3556
rect 28491 3553 28503 3587
rect 28445 3547 28503 3553
rect 30834 3544 30840 3596
rect 30892 3584 30898 3596
rect 31021 3587 31079 3593
rect 31021 3584 31033 3587
rect 30892 3556 31033 3584
rect 30892 3544 30898 3556
rect 31021 3553 31033 3556
rect 31067 3553 31079 3587
rect 31021 3547 31079 3553
rect 32214 3544 32220 3596
rect 32272 3584 32278 3596
rect 33597 3587 33655 3593
rect 33597 3584 33609 3587
rect 32272 3556 33609 3584
rect 32272 3544 32278 3556
rect 33597 3553 33609 3556
rect 33643 3553 33655 3587
rect 33597 3547 33655 3553
rect 33686 3544 33692 3596
rect 33744 3584 33750 3596
rect 36357 3587 36415 3593
rect 36357 3584 36369 3587
rect 33744 3556 36369 3584
rect 33744 3544 33750 3556
rect 36357 3553 36369 3556
rect 36403 3553 36415 3587
rect 36357 3547 36415 3553
rect 38562 3544 38568 3596
rect 38620 3584 38626 3596
rect 39945 3587 40003 3593
rect 39945 3584 39957 3587
rect 38620 3556 39957 3584
rect 38620 3544 38626 3556
rect 39945 3553 39957 3556
rect 39991 3553 40003 3587
rect 39945 3547 40003 3553
rect 41322 3544 41328 3596
rect 41380 3584 41386 3596
rect 42061 3587 42119 3593
rect 42061 3584 42073 3587
rect 41380 3556 42073 3584
rect 41380 3544 41386 3556
rect 42061 3553 42073 3556
rect 42107 3553 42119 3587
rect 42061 3547 42119 3553
rect 10226 3476 10232 3528
rect 10284 3516 10290 3528
rect 10321 3519 10379 3525
rect 10321 3516 10333 3519
rect 10284 3488 10333 3516
rect 10284 3476 10290 3488
rect 10321 3485 10333 3488
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 12158 3476 12164 3528
rect 12216 3516 12222 3528
rect 12253 3519 12311 3525
rect 12253 3516 12265 3519
rect 12216 3488 12265 3516
rect 12216 3476 12222 3488
rect 12253 3485 12265 3488
rect 12299 3485 12311 3519
rect 12253 3479 12311 3485
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 13044 3488 13093 3516
rect 13044 3476 13050 3488
rect 13081 3485 13093 3488
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 14090 3476 14096 3528
rect 14148 3516 14154 3528
rect 14185 3519 14243 3525
rect 14185 3516 14197 3519
rect 14148 3488 14197 3516
rect 14148 3476 14154 3488
rect 14185 3485 14197 3488
rect 14231 3485 14243 3519
rect 14185 3479 14243 3485
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 14976 3488 15025 3516
rect 14976 3476 14982 3488
rect 15013 3485 15025 3488
rect 15059 3485 15071 3519
rect 15013 3479 15071 3485
rect 15746 3476 15752 3528
rect 15804 3516 15810 3528
rect 15841 3519 15899 3525
rect 15841 3516 15853 3519
rect 15804 3488 15853 3516
rect 15804 3476 15810 3488
rect 15841 3485 15853 3488
rect 15887 3485 15899 3519
rect 15841 3479 15899 3485
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 16632 3488 16681 3516
rect 16632 3476 16638 3488
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 17497 3519 17555 3525
rect 17497 3485 17509 3519
rect 17543 3516 17555 3519
rect 17862 3516 17868 3528
rect 17543 3488 17868 3516
rect 17543 3485 17555 3488
rect 17497 3479 17555 3485
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3516 18199 3519
rect 18690 3516 18696 3528
rect 18187 3488 18696 3516
rect 18187 3485 18199 3488
rect 18141 3479 18199 3485
rect 18690 3476 18696 3488
rect 18748 3476 18754 3528
rect 18785 3519 18843 3525
rect 18785 3485 18797 3519
rect 18831 3516 18843 3519
rect 19242 3516 19248 3528
rect 18831 3488 19248 3516
rect 18831 3485 18843 3488
rect 18785 3479 18843 3485
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 20901 3519 20959 3525
rect 20901 3485 20913 3519
rect 20947 3485 20959 3519
rect 20901 3479 20959 3485
rect 21545 3519 21603 3525
rect 21545 3485 21557 3519
rect 21591 3516 21603 3519
rect 22370 3516 22376 3528
rect 21591 3488 22376 3516
rect 21591 3485 21603 3488
rect 21545 3479 21603 3485
rect 20916 3448 20944 3479
rect 22370 3476 22376 3488
rect 22428 3476 22434 3528
rect 30558 3516 30564 3528
rect 30519 3488 30564 3516
rect 30558 3476 30564 3488
rect 30616 3476 30622 3528
rect 33134 3516 33140 3528
rect 33095 3488 33140 3516
rect 33134 3476 33140 3488
rect 33192 3476 33198 3528
rect 35894 3516 35900 3528
rect 35855 3488 35900 3516
rect 35894 3476 35900 3488
rect 35952 3476 35958 3528
rect 39301 3519 39359 3525
rect 39301 3516 39313 3519
rect 37292 3488 39313 3516
rect 24210 3448 24216 3460
rect 20916 3420 24216 3448
rect 24210 3408 24216 3420
rect 24268 3408 24274 3460
rect 24305 3451 24363 3457
rect 24305 3417 24317 3451
rect 24351 3417 24363 3451
rect 25406 3448 25412 3460
rect 25367 3420 25412 3448
rect 24305 3411 24363 3417
rect 22094 3340 22100 3392
rect 22152 3380 22158 3392
rect 23474 3380 23480 3392
rect 22152 3352 23480 3380
rect 22152 3340 22158 3352
rect 23474 3340 23480 3352
rect 23532 3340 23538 3392
rect 24320 3380 24348 3411
rect 25406 3408 25412 3420
rect 25464 3408 25470 3460
rect 27065 3451 27123 3457
rect 27065 3417 27077 3451
rect 27111 3448 27123 3451
rect 28902 3448 28908 3460
rect 27111 3420 28908 3448
rect 27111 3417 27123 3420
rect 27065 3411 27123 3417
rect 28902 3408 28908 3420
rect 28960 3408 28966 3460
rect 30374 3408 30380 3460
rect 30432 3448 30438 3460
rect 30745 3451 30803 3457
rect 30745 3448 30757 3451
rect 30432 3420 30757 3448
rect 30432 3408 30438 3420
rect 30745 3417 30757 3420
rect 30791 3417 30803 3451
rect 30745 3411 30803 3417
rect 33321 3451 33379 3457
rect 33321 3417 33333 3451
rect 33367 3448 33379 3451
rect 33870 3448 33876 3460
rect 33367 3420 33876 3448
rect 33367 3417 33379 3420
rect 33321 3411 33379 3417
rect 33870 3408 33876 3420
rect 33928 3408 33934 3460
rect 36078 3448 36084 3460
rect 36039 3420 36084 3448
rect 36078 3408 36084 3420
rect 36136 3408 36142 3460
rect 36630 3408 36636 3460
rect 36688 3448 36694 3460
rect 37292 3448 37320 3488
rect 39301 3485 39313 3488
rect 39347 3485 39359 3519
rect 39301 3479 39359 3485
rect 40589 3519 40647 3525
rect 40589 3485 40601 3519
rect 40635 3485 40647 3519
rect 40589 3479 40647 3485
rect 42705 3519 42763 3525
rect 42705 3485 42717 3519
rect 42751 3485 42763 3519
rect 42705 3479 42763 3485
rect 36688 3420 37320 3448
rect 36688 3408 36694 3420
rect 38838 3408 38844 3460
rect 38896 3448 38902 3460
rect 40604 3448 40632 3479
rect 38896 3420 40632 3448
rect 38896 3408 38902 3420
rect 41874 3408 41880 3460
rect 41932 3448 41938 3460
rect 42720 3448 42748 3479
rect 43530 3476 43536 3528
rect 43588 3516 43594 3528
rect 44177 3519 44235 3525
rect 44177 3516 44189 3519
rect 43588 3488 44189 3516
rect 43588 3476 43594 3488
rect 44177 3485 44189 3488
rect 44223 3485 44235 3519
rect 44177 3479 44235 3485
rect 44910 3476 44916 3528
rect 44968 3516 44974 3528
rect 45005 3519 45063 3525
rect 45005 3516 45017 3519
rect 44968 3488 45017 3516
rect 44968 3476 44974 3488
rect 45005 3485 45017 3488
rect 45051 3485 45063 3519
rect 45005 3479 45063 3485
rect 46290 3476 46296 3528
rect 46348 3516 46354 3528
rect 46937 3519 46995 3525
rect 46937 3516 46949 3519
rect 46348 3488 46949 3516
rect 46348 3476 46354 3488
rect 46937 3485 46949 3488
rect 46983 3485 46995 3519
rect 46937 3479 46995 3485
rect 47670 3476 47676 3528
rect 47728 3516 47734 3528
rect 47765 3519 47823 3525
rect 47765 3516 47777 3519
rect 47728 3488 47777 3516
rect 47728 3476 47734 3488
rect 47765 3485 47777 3488
rect 47811 3485 47823 3519
rect 47765 3479 47823 3485
rect 49050 3476 49056 3528
rect 49108 3516 49114 3528
rect 49697 3519 49755 3525
rect 49697 3516 49709 3519
rect 49108 3488 49709 3516
rect 49108 3476 49114 3488
rect 49697 3485 49709 3488
rect 49743 3485 49755 3519
rect 49697 3479 49755 3485
rect 50525 3519 50583 3525
rect 50525 3485 50537 3519
rect 50571 3516 50583 3519
rect 50614 3516 50620 3528
rect 50571 3488 50620 3516
rect 50571 3485 50583 3488
rect 50525 3479 50583 3485
rect 50614 3476 50620 3488
rect 50672 3476 50678 3528
rect 51810 3476 51816 3528
rect 51868 3516 51874 3528
rect 52457 3519 52515 3525
rect 52457 3516 52469 3519
rect 51868 3488 52469 3516
rect 51868 3476 51874 3488
rect 52457 3485 52469 3488
rect 52503 3485 52515 3519
rect 52457 3479 52515 3485
rect 41932 3420 42748 3448
rect 41932 3408 41938 3420
rect 26418 3380 26424 3392
rect 24320 3352 26424 3380
rect 26418 3340 26424 3352
rect 26476 3340 26482 3392
rect 35526 3340 35532 3392
rect 35584 3380 35590 3392
rect 40034 3380 40040 3392
rect 35584 3352 40040 3380
rect 35584 3340 35590 3352
rect 40034 3340 40040 3352
rect 40092 3340 40098 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 22186 3176 22192 3188
rect 22147 3148 22192 3176
rect 22186 3136 22192 3148
rect 22244 3136 22250 3188
rect 24486 3176 24492 3188
rect 23308 3148 24492 3176
rect 23308 3108 23336 3148
rect 24486 3136 24492 3148
rect 24544 3136 24550 3188
rect 33042 3136 33048 3188
rect 33100 3176 33106 3188
rect 33594 3176 33600 3188
rect 33100 3148 33600 3176
rect 33100 3136 33106 3148
rect 33594 3136 33600 3148
rect 33652 3136 33658 3188
rect 35342 3136 35348 3188
rect 35400 3176 35406 3188
rect 39298 3176 39304 3188
rect 35400 3148 39304 3176
rect 35400 3136 35406 3148
rect 39298 3136 39304 3148
rect 39356 3136 39362 3188
rect 24026 3108 24032 3120
rect 20180 3080 23336 3108
rect 23987 3080 24032 3108
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2972 17463 2975
rect 18966 2972 18972 2984
rect 17451 2944 18972 2972
rect 17451 2941 17463 2944
rect 17405 2935 17463 2941
rect 18966 2932 18972 2944
rect 19024 2932 19030 2984
rect 20180 2981 20208 3080
rect 24026 3068 24032 3080
rect 24084 3068 24090 3120
rect 25685 3111 25743 3117
rect 25685 3077 25697 3111
rect 25731 3108 25743 3111
rect 27246 3108 27252 3120
rect 25731 3080 27252 3108
rect 25731 3077 25743 3080
rect 25685 3071 25743 3077
rect 27246 3068 27252 3080
rect 27304 3068 27310 3120
rect 34146 3068 34152 3120
rect 34204 3108 34210 3120
rect 34204 3080 35940 3108
rect 34204 3068 34210 3080
rect 21637 3043 21695 3049
rect 21637 3009 21649 3043
rect 21683 3040 21695 3043
rect 22094 3040 22100 3052
rect 21683 3012 22100 3040
rect 21683 3009 21695 3012
rect 21637 3003 21695 3009
rect 22094 3000 22100 3012
rect 22152 3040 22158 3052
rect 22152 3012 22197 3040
rect 22152 3000 22158 3012
rect 22370 3000 22376 3052
rect 22428 3040 22434 3052
rect 23845 3043 23903 3049
rect 23845 3040 23857 3043
rect 22428 3012 23857 3040
rect 22428 3000 22434 3012
rect 23845 3009 23857 3012
rect 23891 3009 23903 3043
rect 23845 3003 23903 3009
rect 20165 2975 20223 2981
rect 20165 2941 20177 2975
rect 20211 2941 20223 2975
rect 20165 2935 20223 2941
rect 20993 2975 21051 2981
rect 20993 2941 21005 2975
rect 21039 2972 21051 2975
rect 25038 2972 25044 2984
rect 21039 2944 25044 2972
rect 21039 2941 21051 2944
rect 20993 2935 21051 2941
rect 25038 2932 25044 2944
rect 25096 2932 25102 2984
rect 26602 2972 26608 2984
rect 26563 2944 26608 2972
rect 26602 2932 26608 2944
rect 26660 2932 26666 2984
rect 26786 2972 26792 2984
rect 26747 2944 26792 2972
rect 26786 2932 26792 2944
rect 26844 2932 26850 2984
rect 28445 2975 28503 2981
rect 28445 2941 28457 2975
rect 28491 2941 28503 2975
rect 28445 2935 28503 2941
rect 18233 2907 18291 2913
rect 18233 2873 18245 2907
rect 18279 2904 18291 2907
rect 19426 2904 19432 2916
rect 18279 2876 19432 2904
rect 18279 2873 18291 2876
rect 18233 2867 18291 2873
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 19521 2907 19579 2913
rect 19521 2873 19533 2907
rect 19567 2904 19579 2907
rect 22738 2904 22744 2916
rect 19567 2876 22744 2904
rect 19567 2873 19579 2876
rect 19521 2867 19579 2873
rect 22738 2864 22744 2876
rect 22796 2864 22802 2916
rect 25498 2904 25504 2916
rect 22848 2876 25504 2904
rect 8481 2839 8539 2845
rect 8481 2805 8493 2839
rect 8527 2836 8539 2839
rect 8570 2836 8576 2848
rect 8527 2808 8576 2836
rect 8527 2805 8539 2808
rect 8481 2799 8539 2805
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 9125 2839 9183 2845
rect 9125 2805 9137 2839
rect 9171 2836 9183 2839
rect 9306 2836 9312 2848
rect 9171 2808 9312 2836
rect 9171 2805 9183 2808
rect 9125 2799 9183 2805
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 9950 2836 9956 2848
rect 9911 2808 9956 2836
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 10597 2839 10655 2845
rect 10597 2805 10609 2839
rect 10643 2836 10655 2839
rect 10778 2836 10784 2848
rect 10643 2808 10784 2836
rect 10643 2805 10655 2808
rect 10597 2799 10655 2805
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 11241 2839 11299 2845
rect 11241 2805 11253 2839
rect 11287 2836 11299 2839
rect 11330 2836 11336 2848
rect 11287 2808 11336 2836
rect 11287 2805 11299 2808
rect 11241 2799 11299 2805
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 11701 2839 11759 2845
rect 11701 2836 11713 2839
rect 11664 2808 11713 2836
rect 11664 2796 11670 2808
rect 11701 2805 11713 2808
rect 11747 2805 11759 2839
rect 12710 2836 12716 2848
rect 12671 2808 12716 2836
rect 11701 2799 11759 2805
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 13357 2839 13415 2845
rect 13357 2805 13369 2839
rect 13403 2836 13415 2839
rect 13538 2836 13544 2848
rect 13403 2808 13544 2836
rect 13403 2805 13415 2808
rect 13357 2799 13415 2805
rect 13538 2796 13544 2808
rect 13596 2796 13602 2848
rect 14001 2839 14059 2845
rect 14001 2805 14013 2839
rect 14047 2836 14059 2839
rect 14366 2836 14372 2848
rect 14047 2808 14372 2836
rect 14047 2805 14059 2808
rect 14001 2799 14059 2805
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 14645 2839 14703 2845
rect 14645 2805 14657 2839
rect 14691 2836 14703 2839
rect 15194 2836 15200 2848
rect 14691 2808 15200 2836
rect 14691 2805 14703 2808
rect 14645 2799 14703 2805
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 15473 2839 15531 2845
rect 15473 2805 15485 2839
rect 15519 2836 15531 2839
rect 16022 2836 16028 2848
rect 15519 2808 16028 2836
rect 15519 2805 15531 2808
rect 15473 2799 15531 2805
rect 16022 2796 16028 2808
rect 16080 2796 16086 2848
rect 16117 2839 16175 2845
rect 16117 2805 16129 2839
rect 16163 2836 16175 2839
rect 16298 2836 16304 2848
rect 16163 2808 16304 2836
rect 16163 2805 16175 2808
rect 16117 2799 16175 2805
rect 16298 2796 16304 2808
rect 16356 2796 16362 2848
rect 16761 2839 16819 2845
rect 16761 2805 16773 2839
rect 16807 2836 16819 2839
rect 17310 2836 17316 2848
rect 16807 2808 17316 2836
rect 16807 2805 16819 2808
rect 16761 2799 16819 2805
rect 17310 2796 17316 2808
rect 17368 2796 17374 2848
rect 18877 2839 18935 2845
rect 18877 2805 18889 2839
rect 18923 2836 18935 2839
rect 20898 2836 20904 2848
rect 18923 2808 20904 2836
rect 18923 2805 18935 2808
rect 18877 2799 18935 2805
rect 20898 2796 20904 2808
rect 20956 2796 20962 2848
rect 21545 2839 21603 2845
rect 21545 2805 21557 2839
rect 21591 2836 21603 2839
rect 22848 2836 22876 2876
rect 25498 2864 25504 2876
rect 25556 2864 25562 2916
rect 28460 2904 28488 2935
rect 28534 2932 28540 2984
rect 28592 2972 28598 2984
rect 29365 2975 29423 2981
rect 29365 2972 29377 2975
rect 28592 2944 29377 2972
rect 28592 2932 28598 2944
rect 29365 2941 29377 2944
rect 29411 2941 29423 2975
rect 29546 2972 29552 2984
rect 29507 2944 29552 2972
rect 29365 2935 29423 2941
rect 29546 2932 29552 2944
rect 29604 2932 29610 2984
rect 31110 2972 31116 2984
rect 31071 2944 31116 2972
rect 31110 2932 31116 2944
rect 31168 2932 31174 2984
rect 31938 2972 31944 2984
rect 31899 2944 31944 2972
rect 31938 2932 31944 2944
rect 31996 2932 32002 2984
rect 33410 2972 33416 2984
rect 33371 2944 33416 2972
rect 33410 2932 33416 2944
rect 33468 2932 33474 2984
rect 33594 2972 33600 2984
rect 33555 2944 33600 2972
rect 33594 2932 33600 2944
rect 33652 2932 33658 2984
rect 34514 2972 34520 2984
rect 34475 2944 34520 2972
rect 34514 2932 34520 2944
rect 34572 2932 34578 2984
rect 34698 2972 34704 2984
rect 34659 2944 34704 2972
rect 34698 2932 34704 2944
rect 34756 2932 34762 2984
rect 34977 2975 35035 2981
rect 34977 2941 34989 2975
rect 35023 2941 35035 2975
rect 34977 2935 35035 2941
rect 29454 2904 29460 2916
rect 28460 2876 29460 2904
rect 29454 2864 29460 2876
rect 29512 2864 29518 2916
rect 32490 2864 32496 2916
rect 32548 2904 32554 2916
rect 34992 2904 35020 2935
rect 32548 2876 35020 2904
rect 35912 2904 35940 3080
rect 36354 3068 36360 3120
rect 36412 3108 36418 3120
rect 36412 3080 39252 3108
rect 36412 3068 36418 3080
rect 37274 3040 37280 3052
rect 37235 3012 37280 3040
rect 37274 3000 37280 3012
rect 37332 3000 37338 3052
rect 37458 2972 37464 2984
rect 37419 2944 37464 2972
rect 37458 2932 37464 2944
rect 37516 2932 37522 2984
rect 37737 2975 37795 2981
rect 37737 2941 37749 2975
rect 37783 2941 37795 2975
rect 39224 2972 39252 3080
rect 39666 3000 39672 3052
rect 39724 3040 39730 3052
rect 41325 3043 41383 3049
rect 41325 3040 41337 3043
rect 39724 3012 41337 3040
rect 39724 3000 39730 3012
rect 41325 3009 41337 3012
rect 41371 3009 41383 3043
rect 41325 3003 41383 3009
rect 40037 2975 40095 2981
rect 40037 2972 40049 2975
rect 39224 2944 40049 2972
rect 37737 2935 37795 2941
rect 40037 2941 40049 2944
rect 40083 2941 40095 2975
rect 40037 2935 40095 2941
rect 37752 2904 37780 2935
rect 40218 2932 40224 2984
rect 40276 2972 40282 2984
rect 41969 2975 42027 2981
rect 41969 2972 41981 2975
rect 40276 2944 41981 2972
rect 40276 2932 40282 2944
rect 41969 2941 41981 2944
rect 42015 2941 42027 2975
rect 41969 2935 42027 2941
rect 42150 2932 42156 2984
rect 42208 2972 42214 2984
rect 43441 2975 43499 2981
rect 43441 2972 43453 2975
rect 42208 2944 43453 2972
rect 42208 2932 42214 2944
rect 43441 2941 43453 2944
rect 43487 2941 43499 2975
rect 43441 2935 43499 2941
rect 44634 2932 44640 2984
rect 44692 2972 44698 2984
rect 45557 2975 45615 2981
rect 45557 2972 45569 2975
rect 44692 2944 45569 2972
rect 44692 2932 44698 2944
rect 45557 2941 45569 2944
rect 45603 2941 45615 2975
rect 45557 2935 45615 2941
rect 35912 2876 37780 2904
rect 32548 2864 32554 2876
rect 38010 2864 38016 2916
rect 38068 2904 38074 2916
rect 40681 2907 40739 2913
rect 40681 2904 40693 2907
rect 38068 2876 40693 2904
rect 38068 2864 38074 2876
rect 40681 2873 40693 2876
rect 40727 2873 40739 2907
rect 40681 2867 40739 2873
rect 41046 2864 41052 2916
rect 41104 2904 41110 2916
rect 41104 2876 41414 2904
rect 41104 2864 41110 2876
rect 21591 2808 22876 2836
rect 22925 2839 22983 2845
rect 21591 2805 21603 2808
rect 21545 2799 21603 2805
rect 22925 2805 22937 2839
rect 22971 2836 22983 2839
rect 27890 2836 27896 2848
rect 22971 2808 27896 2836
rect 22971 2805 22983 2808
rect 22925 2799 22983 2805
rect 27890 2796 27896 2808
rect 27948 2796 27954 2848
rect 31386 2796 31392 2848
rect 31444 2836 31450 2848
rect 31754 2836 31760 2848
rect 31444 2808 31760 2836
rect 31444 2796 31450 2808
rect 31754 2796 31760 2808
rect 31812 2796 31818 2848
rect 34790 2796 34796 2848
rect 34848 2836 34854 2848
rect 38654 2836 38660 2848
rect 34848 2808 38660 2836
rect 34848 2796 34854 2808
rect 38654 2796 38660 2808
rect 38712 2796 38718 2848
rect 41386 2836 41414 2876
rect 43254 2864 43260 2916
rect 43312 2904 43318 2916
rect 44085 2907 44143 2913
rect 44085 2904 44097 2907
rect 43312 2876 44097 2904
rect 43312 2864 43318 2876
rect 44085 2873 44097 2876
rect 44131 2873 44143 2907
rect 44085 2867 44143 2873
rect 45462 2864 45468 2916
rect 45520 2904 45526 2916
rect 46201 2907 46259 2913
rect 46201 2904 46213 2907
rect 45520 2876 46213 2904
rect 45520 2864 45526 2876
rect 46201 2873 46213 2876
rect 46247 2873 46259 2907
rect 46201 2867 46259 2873
rect 46566 2864 46572 2916
rect 46624 2904 46630 2916
rect 47489 2907 47547 2913
rect 47489 2904 47501 2907
rect 46624 2876 47501 2904
rect 46624 2864 46630 2876
rect 47489 2873 47501 2876
rect 47535 2873 47547 2907
rect 47489 2867 47547 2873
rect 48222 2864 48228 2916
rect 48280 2904 48286 2916
rect 48961 2907 49019 2913
rect 48961 2904 48973 2907
rect 48280 2876 48973 2904
rect 48280 2864 48286 2876
rect 48961 2873 48973 2876
rect 49007 2873 49019 2907
rect 48961 2867 49019 2873
rect 49326 2864 49332 2916
rect 49384 2904 49390 2916
rect 50249 2907 50307 2913
rect 50249 2904 50261 2907
rect 49384 2876 50261 2904
rect 49384 2864 49390 2876
rect 50249 2873 50261 2876
rect 50295 2873 50307 2907
rect 50249 2867 50307 2873
rect 50982 2864 50988 2916
rect 51040 2904 51046 2916
rect 51721 2907 51779 2913
rect 51721 2904 51733 2907
rect 51040 2876 51733 2904
rect 51040 2864 51046 2876
rect 51721 2873 51733 2876
rect 51767 2873 51779 2907
rect 51721 2867 51779 2873
rect 52086 2864 52092 2916
rect 52144 2904 52150 2916
rect 53009 2907 53067 2913
rect 53009 2904 53021 2907
rect 52144 2876 53021 2904
rect 52144 2864 52150 2876
rect 53009 2873 53021 2876
rect 53055 2873 53067 2907
rect 53009 2867 53067 2873
rect 42797 2839 42855 2845
rect 42797 2836 42809 2839
rect 41386 2808 42809 2836
rect 42797 2805 42809 2808
rect 42843 2805 42855 2839
rect 42797 2799 42855 2805
rect 43806 2796 43812 2848
rect 43864 2836 43870 2848
rect 44729 2839 44787 2845
rect 44729 2836 44741 2839
rect 43864 2808 44741 2836
rect 43864 2796 43870 2808
rect 44729 2805 44741 2808
rect 44775 2805 44787 2839
rect 44729 2799 44787 2805
rect 46014 2796 46020 2848
rect 46072 2836 46078 2848
rect 46845 2839 46903 2845
rect 46845 2836 46857 2839
rect 46072 2808 46857 2836
rect 46072 2796 46078 2808
rect 46845 2805 46857 2808
rect 46891 2805 46903 2839
rect 46845 2799 46903 2805
rect 47394 2796 47400 2848
rect 47452 2836 47458 2848
rect 48317 2839 48375 2845
rect 48317 2836 48329 2839
rect 47452 2808 48329 2836
rect 47452 2796 47458 2808
rect 48317 2805 48329 2808
rect 48363 2805 48375 2839
rect 48317 2799 48375 2805
rect 48774 2796 48780 2848
rect 48832 2836 48838 2848
rect 49605 2839 49663 2845
rect 49605 2836 49617 2839
rect 48832 2808 49617 2836
rect 48832 2796 48838 2808
rect 49605 2805 49617 2808
rect 49651 2805 49663 2839
rect 49605 2799 49663 2805
rect 50154 2796 50160 2848
rect 50212 2836 50218 2848
rect 51077 2839 51135 2845
rect 51077 2836 51089 2839
rect 50212 2808 51089 2836
rect 50212 2796 50218 2808
rect 51077 2805 51089 2808
rect 51123 2805 51135 2839
rect 51077 2799 51135 2805
rect 51534 2796 51540 2848
rect 51592 2836 51598 2848
rect 52365 2839 52423 2845
rect 52365 2836 52377 2839
rect 51592 2808 52377 2836
rect 51592 2796 51598 2808
rect 52365 2805 52377 2808
rect 52411 2805 52423 2839
rect 52365 2799 52423 2805
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 16761 2635 16819 2641
rect 16761 2601 16773 2635
rect 16807 2632 16819 2635
rect 18138 2632 18144 2644
rect 16807 2604 18144 2632
rect 16807 2601 16819 2604
rect 16761 2595 16819 2601
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 22281 2635 22339 2641
rect 22281 2601 22293 2635
rect 22327 2632 22339 2635
rect 22738 2632 22744 2644
rect 22327 2604 22744 2632
rect 22327 2601 22339 2604
rect 22281 2595 22339 2601
rect 22738 2592 22744 2604
rect 22796 2592 22802 2644
rect 22925 2635 22983 2641
rect 22925 2601 22937 2635
rect 22971 2632 22983 2635
rect 23842 2632 23848 2644
rect 22971 2604 23848 2632
rect 22971 2601 22983 2604
rect 22925 2595 22983 2601
rect 23842 2592 23848 2604
rect 23900 2592 23906 2644
rect 24305 2635 24363 2641
rect 24305 2601 24317 2635
rect 24351 2632 24363 2635
rect 25314 2632 25320 2644
rect 24351 2604 25320 2632
rect 24351 2601 24363 2604
rect 24305 2595 24363 2601
rect 25314 2592 25320 2604
rect 25372 2592 25378 2644
rect 25685 2635 25743 2641
rect 25685 2601 25697 2635
rect 25731 2632 25743 2635
rect 26602 2632 26608 2644
rect 25731 2604 26608 2632
rect 25731 2601 25743 2604
rect 25685 2595 25743 2601
rect 26602 2592 26608 2604
rect 26660 2592 26666 2644
rect 27065 2635 27123 2641
rect 27065 2601 27077 2635
rect 27111 2632 27123 2635
rect 28534 2632 28540 2644
rect 27111 2604 28540 2632
rect 27111 2601 27123 2604
rect 27065 2595 27123 2601
rect 28534 2592 28540 2604
rect 28592 2592 28598 2644
rect 29733 2635 29791 2641
rect 29733 2601 29745 2635
rect 29779 2632 29791 2635
rect 30374 2632 30380 2644
rect 29779 2604 30380 2632
rect 29779 2601 29791 2604
rect 29733 2595 29791 2601
rect 30374 2592 30380 2604
rect 30432 2592 30438 2644
rect 30558 2592 30564 2644
rect 30616 2632 30622 2644
rect 30653 2635 30711 2641
rect 30653 2632 30665 2635
rect 30616 2604 30665 2632
rect 30616 2592 30622 2604
rect 30653 2601 30665 2604
rect 30699 2601 30711 2635
rect 30653 2595 30711 2601
rect 32585 2635 32643 2641
rect 32585 2601 32597 2635
rect 32631 2632 32643 2635
rect 33134 2632 33140 2644
rect 32631 2604 33140 2632
rect 32631 2601 32643 2604
rect 32585 2595 32643 2601
rect 33134 2592 33140 2604
rect 33192 2592 33198 2644
rect 33229 2635 33287 2641
rect 33229 2601 33241 2635
rect 33275 2632 33287 2635
rect 33410 2632 33416 2644
rect 33275 2604 33416 2632
rect 33275 2601 33287 2604
rect 33229 2595 33287 2601
rect 33410 2592 33416 2604
rect 33468 2592 33474 2644
rect 33870 2632 33876 2644
rect 33831 2604 33876 2632
rect 33870 2592 33876 2604
rect 33928 2592 33934 2644
rect 34514 2632 34520 2644
rect 34475 2604 34520 2632
rect 34514 2592 34520 2604
rect 34572 2592 34578 2644
rect 34698 2592 34704 2644
rect 34756 2632 34762 2644
rect 35253 2635 35311 2641
rect 35253 2632 35265 2635
rect 34756 2604 35265 2632
rect 34756 2592 34762 2604
rect 35253 2601 35265 2604
rect 35299 2601 35311 2635
rect 35253 2595 35311 2601
rect 35989 2635 36047 2641
rect 35989 2601 36001 2635
rect 36035 2632 36047 2635
rect 36078 2632 36084 2644
rect 36035 2604 36084 2632
rect 36035 2601 36047 2604
rect 35989 2595 36047 2601
rect 36078 2592 36084 2604
rect 36136 2592 36142 2644
rect 37369 2635 37427 2641
rect 37369 2601 37381 2635
rect 37415 2632 37427 2635
rect 37458 2632 37464 2644
rect 37415 2604 37464 2632
rect 37415 2601 37427 2604
rect 37369 2595 37427 2601
rect 37458 2592 37464 2604
rect 37516 2592 37522 2644
rect 37918 2592 37924 2644
rect 37976 2632 37982 2644
rect 38013 2635 38071 2641
rect 38013 2632 38025 2635
rect 37976 2604 38025 2632
rect 37976 2592 37982 2604
rect 38013 2601 38025 2604
rect 38059 2601 38071 2635
rect 38654 2632 38660 2644
rect 38615 2604 38660 2632
rect 38013 2595 38071 2601
rect 38654 2592 38660 2604
rect 38712 2592 38718 2644
rect 39298 2632 39304 2644
rect 39259 2604 39304 2632
rect 39298 2592 39304 2604
rect 39356 2592 39362 2644
rect 40034 2632 40040 2644
rect 39995 2604 40040 2632
rect 40034 2592 40040 2604
rect 40092 2592 40098 2644
rect 47118 2592 47124 2644
rect 47176 2632 47182 2644
rect 48961 2635 49019 2641
rect 48961 2632 48973 2635
rect 47176 2604 48973 2632
rect 47176 2592 47182 2604
rect 48961 2601 48973 2604
rect 49007 2601 49019 2635
rect 48961 2595 49019 2601
rect 49878 2592 49884 2644
rect 49936 2632 49942 2644
rect 51721 2635 51779 2641
rect 51721 2632 51733 2635
rect 49936 2604 51733 2632
rect 49936 2592 49942 2604
rect 51721 2601 51733 2604
rect 51767 2601 51779 2635
rect 51721 2595 51779 2601
rect 9861 2567 9919 2573
rect 9861 2533 9873 2567
rect 9907 2564 9919 2567
rect 10502 2564 10508 2576
rect 9907 2536 10508 2564
rect 9907 2533 9919 2536
rect 9861 2527 9919 2533
rect 10502 2524 10508 2536
rect 10560 2524 10566 2576
rect 11241 2567 11299 2573
rect 11241 2533 11253 2567
rect 11287 2564 11299 2567
rect 11882 2564 11888 2576
rect 11287 2536 11888 2564
rect 11287 2533 11299 2536
rect 11241 2527 11299 2533
rect 11882 2524 11888 2536
rect 11940 2524 11946 2576
rect 12621 2567 12679 2573
rect 12621 2533 12633 2567
rect 12667 2564 12679 2567
rect 13262 2564 13268 2576
rect 12667 2536 13268 2564
rect 12667 2533 12679 2536
rect 12621 2527 12679 2533
rect 13262 2524 13268 2536
rect 13320 2524 13326 2576
rect 14001 2567 14059 2573
rect 14001 2533 14013 2567
rect 14047 2564 14059 2567
rect 14642 2564 14648 2576
rect 14047 2536 14648 2564
rect 14047 2533 14059 2536
rect 14001 2527 14059 2533
rect 14642 2524 14648 2536
rect 14700 2524 14706 2576
rect 16025 2567 16083 2573
rect 16025 2533 16037 2567
rect 16071 2564 16083 2567
rect 17586 2564 17592 2576
rect 16071 2536 17592 2564
rect 16071 2533 16083 2536
rect 16025 2527 16083 2533
rect 17586 2524 17592 2536
rect 17644 2524 17650 2576
rect 18785 2567 18843 2573
rect 18785 2533 18797 2567
rect 18831 2564 18843 2567
rect 23106 2564 23112 2576
rect 18831 2536 23112 2564
rect 18831 2533 18843 2536
rect 18785 2527 18843 2533
rect 23106 2524 23112 2536
rect 23164 2524 23170 2576
rect 23569 2567 23627 2573
rect 23569 2533 23581 2567
rect 23615 2564 23627 2567
rect 25406 2564 25412 2576
rect 23615 2536 25412 2564
rect 23615 2533 23627 2536
rect 23569 2527 23627 2533
rect 25406 2524 25412 2536
rect 25464 2524 25470 2576
rect 26329 2567 26387 2573
rect 26329 2533 26341 2567
rect 26375 2564 26387 2567
rect 26786 2564 26792 2576
rect 26375 2536 26792 2564
rect 26375 2533 26387 2536
rect 26329 2527 26387 2533
rect 26786 2524 26792 2536
rect 26844 2524 26850 2576
rect 27709 2567 27767 2573
rect 27709 2533 27721 2567
rect 27755 2564 27767 2567
rect 29546 2564 29552 2576
rect 27755 2536 29552 2564
rect 27755 2533 27767 2536
rect 27709 2527 27767 2533
rect 29546 2524 29552 2536
rect 29604 2524 29610 2576
rect 31941 2567 31999 2573
rect 31941 2533 31953 2567
rect 31987 2564 31999 2567
rect 33594 2564 33600 2576
rect 31987 2536 33600 2564
rect 31987 2533 31999 2536
rect 31941 2527 31999 2533
rect 33594 2524 33600 2536
rect 33652 2524 33658 2576
rect 35894 2524 35900 2576
rect 35952 2564 35958 2576
rect 36541 2567 36599 2573
rect 36541 2564 36553 2567
rect 35952 2536 36553 2564
rect 35952 2524 35958 2536
rect 36541 2533 36553 2536
rect 36587 2533 36599 2567
rect 36541 2527 36599 2533
rect 39390 2524 39396 2576
rect 39448 2564 39454 2576
rect 42061 2567 42119 2573
rect 42061 2564 42073 2567
rect 39448 2536 42073 2564
rect 39448 2524 39454 2536
rect 42061 2533 42073 2536
rect 42107 2533 42119 2567
rect 42061 2527 42119 2533
rect 42426 2524 42432 2576
rect 42484 2564 42490 2576
rect 44177 2567 44235 2573
rect 44177 2564 44189 2567
rect 42484 2536 44189 2564
rect 42484 2524 42490 2536
rect 44177 2533 44189 2536
rect 44223 2533 44235 2567
rect 44177 2527 44235 2533
rect 45186 2524 45192 2576
rect 45244 2564 45250 2576
rect 46937 2567 46995 2573
rect 46937 2564 46949 2567
rect 45244 2536 46949 2564
rect 45244 2524 45250 2536
rect 46937 2533 46949 2536
rect 46983 2533 46995 2567
rect 46937 2527 46995 2533
rect 47946 2524 47952 2576
rect 48004 2564 48010 2576
rect 49697 2567 49755 2573
rect 49697 2564 49709 2567
rect 48004 2536 49709 2564
rect 48004 2524 48010 2536
rect 49697 2533 49709 2536
rect 49743 2533 49755 2567
rect 49697 2527 49755 2533
rect 51258 2524 51264 2576
rect 51316 2564 51322 2576
rect 53101 2567 53159 2573
rect 53101 2564 53113 2567
rect 51316 2536 53113 2564
rect 51316 2524 51322 2536
rect 53101 2533 53113 2536
rect 53147 2533 53159 2567
rect 53101 2527 53159 2533
rect 15381 2499 15439 2505
rect 15381 2465 15393 2499
rect 15427 2496 15439 2499
rect 16850 2496 16856 2508
rect 15427 2468 16856 2496
rect 15427 2465 15439 2468
rect 15381 2459 15439 2465
rect 16850 2456 16856 2468
rect 16908 2456 16914 2508
rect 17405 2499 17463 2505
rect 17405 2465 17417 2499
rect 17451 2496 17463 2499
rect 19334 2496 19340 2508
rect 17451 2468 19340 2496
rect 17451 2465 17463 2468
rect 17405 2459 17463 2465
rect 19334 2456 19340 2468
rect 19392 2456 19398 2508
rect 20165 2499 20223 2505
rect 20165 2465 20177 2499
rect 20211 2496 20223 2499
rect 21545 2499 21603 2505
rect 20211 2468 21496 2496
rect 20211 2465 20223 2468
rect 20165 2459 20223 2465
rect 7101 2431 7159 2437
rect 7101 2397 7113 2431
rect 7147 2428 7159 2431
rect 7650 2428 7656 2440
rect 7147 2400 7656 2428
rect 7147 2397 7159 2400
rect 7101 2391 7159 2397
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2428 7803 2431
rect 8202 2428 8208 2440
rect 7791 2400 8208 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2428 8539 2431
rect 8938 2428 8944 2440
rect 8527 2400 8944 2428
rect 8527 2397 8539 2400
rect 8481 2391 8539 2397
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9674 2428 9680 2440
rect 9171 2400 9680 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 11054 2428 11060 2440
rect 10551 2400 11060 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2428 11943 2431
rect 12434 2428 12440 2440
rect 11931 2400 12440 2428
rect 11931 2397 11943 2400
rect 11885 2391 11943 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2428 13323 2431
rect 13814 2428 13820 2440
rect 13311 2400 13820 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 13814 2388 13820 2400
rect 13872 2388 13878 2440
rect 14645 2431 14703 2437
rect 14645 2397 14657 2431
rect 14691 2428 14703 2431
rect 15470 2428 15476 2440
rect 14691 2400 15476 2428
rect 14691 2397 14703 2400
rect 14645 2391 14703 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 18141 2431 18199 2437
rect 18141 2397 18153 2431
rect 18187 2397 18199 2431
rect 18141 2391 18199 2397
rect 19521 2431 19579 2437
rect 19521 2397 19533 2431
rect 19567 2428 19579 2431
rect 19978 2428 19984 2440
rect 19567 2400 19984 2428
rect 19567 2397 19579 2400
rect 19521 2391 19579 2397
rect 18156 2360 18184 2391
rect 19978 2388 19984 2400
rect 20036 2388 20042 2440
rect 20901 2431 20959 2437
rect 20901 2397 20913 2431
rect 20947 2428 20959 2431
rect 21358 2428 21364 2440
rect 20947 2400 21364 2428
rect 20947 2397 20959 2400
rect 20901 2391 20959 2397
rect 21358 2388 21364 2400
rect 21416 2388 21422 2440
rect 21468 2428 21496 2468
rect 21545 2465 21557 2499
rect 21591 2496 21603 2499
rect 24854 2496 24860 2508
rect 21591 2468 24860 2496
rect 21591 2465 21603 2468
rect 21545 2459 21603 2465
rect 24854 2456 24860 2468
rect 24912 2456 24918 2508
rect 24949 2499 25007 2505
rect 24949 2465 24961 2499
rect 24995 2496 25007 2499
rect 26510 2496 26516 2508
rect 24995 2468 26516 2496
rect 24995 2465 25007 2468
rect 24949 2459 25007 2465
rect 26510 2456 26516 2468
rect 26568 2456 26574 2508
rect 29181 2499 29239 2505
rect 29181 2465 29193 2499
rect 29227 2496 29239 2499
rect 30466 2496 30472 2508
rect 29227 2468 30472 2496
rect 29227 2465 29239 2468
rect 29181 2459 29239 2465
rect 30466 2456 30472 2468
rect 30524 2456 30530 2508
rect 37182 2456 37188 2508
rect 37240 2496 37246 2508
rect 40681 2499 40739 2505
rect 40681 2496 40693 2499
rect 37240 2468 40693 2496
rect 37240 2456 37246 2468
rect 40681 2465 40693 2468
rect 40727 2465 40739 2499
rect 40681 2459 40739 2465
rect 41598 2456 41604 2508
rect 41656 2496 41662 2508
rect 43441 2499 43499 2505
rect 43441 2496 43453 2499
rect 41656 2468 43453 2496
rect 41656 2456 41662 2468
rect 43441 2465 43453 2468
rect 43487 2465 43499 2499
rect 43441 2459 43499 2465
rect 44082 2456 44088 2508
rect 44140 2496 44146 2508
rect 45557 2499 45615 2505
rect 45557 2496 45569 2499
rect 44140 2468 45569 2496
rect 44140 2456 44146 2468
rect 45557 2465 45569 2468
rect 45603 2465 45615 2499
rect 45557 2459 45615 2465
rect 46842 2456 46848 2508
rect 46900 2496 46906 2508
rect 48317 2499 48375 2505
rect 48317 2496 48329 2499
rect 46900 2468 48329 2496
rect 46900 2456 46906 2468
rect 48317 2465 48329 2468
rect 48363 2465 48375 2499
rect 48317 2459 48375 2465
rect 49602 2456 49608 2508
rect 49660 2496 49666 2508
rect 51077 2499 51135 2505
rect 51077 2496 51089 2499
rect 49660 2468 51089 2496
rect 49660 2456 49666 2468
rect 51077 2465 51089 2468
rect 51123 2465 51135 2499
rect 51077 2459 51135 2465
rect 52362 2456 52368 2508
rect 52420 2496 52426 2508
rect 53837 2499 53895 2505
rect 53837 2496 53849 2499
rect 52420 2468 53849 2496
rect 52420 2456 52426 2468
rect 53837 2465 53849 2468
rect 53883 2465 53895 2499
rect 53837 2459 53895 2465
rect 21468 2400 23428 2428
rect 21450 2360 21456 2372
rect 18156 2332 21456 2360
rect 21450 2320 21456 2332
rect 21508 2320 21514 2372
rect 23400 2360 23428 2400
rect 23474 2388 23480 2440
rect 23532 2428 23538 2440
rect 25041 2431 25099 2437
rect 23532 2400 23577 2428
rect 23532 2388 23538 2400
rect 25041 2397 25053 2431
rect 25087 2428 25099 2431
rect 26237 2431 26295 2437
rect 26237 2428 26249 2431
rect 25087 2400 26249 2428
rect 25087 2397 25099 2400
rect 25041 2391 25099 2397
rect 26237 2397 26249 2400
rect 26283 2428 26295 2431
rect 27617 2431 27675 2437
rect 27617 2428 27629 2431
rect 26283 2400 27629 2428
rect 26283 2397 26295 2400
rect 26237 2391 26295 2397
rect 27617 2397 27629 2400
rect 27663 2428 27675 2431
rect 28261 2431 28319 2437
rect 28261 2428 28273 2431
rect 27663 2400 28273 2428
rect 27663 2397 27675 2400
rect 27617 2391 27675 2397
rect 28261 2397 28273 2400
rect 28307 2428 28319 2431
rect 29638 2428 29644 2440
rect 28307 2400 29644 2428
rect 28307 2397 28319 2400
rect 28261 2391 28319 2397
rect 29638 2388 29644 2400
rect 29696 2388 29702 2440
rect 32950 2388 32956 2440
rect 33008 2428 33014 2440
rect 33321 2431 33379 2437
rect 33321 2428 33333 2431
rect 33008 2400 33333 2428
rect 33008 2388 33014 2400
rect 33321 2397 33333 2400
rect 33367 2428 33379 2431
rect 33965 2431 34023 2437
rect 33965 2428 33977 2431
rect 33367 2400 33977 2428
rect 33367 2397 33379 2400
rect 33321 2391 33379 2397
rect 33965 2397 33977 2400
rect 34011 2428 34023 2431
rect 35345 2431 35403 2437
rect 35345 2428 35357 2431
rect 34011 2400 35357 2428
rect 34011 2397 34023 2400
rect 33965 2391 34023 2397
rect 35345 2397 35357 2400
rect 35391 2428 35403 2431
rect 35897 2431 35955 2437
rect 35897 2428 35909 2431
rect 35391 2400 35909 2428
rect 35391 2397 35403 2400
rect 35345 2391 35403 2397
rect 35897 2397 35909 2400
rect 35943 2428 35955 2431
rect 36722 2428 36728 2440
rect 35943 2400 36728 2428
rect 35943 2397 35955 2400
rect 35897 2391 35955 2397
rect 36722 2388 36728 2400
rect 36780 2428 36786 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36780 2400 37289 2428
rect 36780 2388 36786 2400
rect 37277 2397 37289 2400
rect 37323 2428 37335 2431
rect 37921 2431 37979 2437
rect 37921 2428 37933 2431
rect 37323 2400 37933 2428
rect 37323 2397 37335 2400
rect 37277 2391 37335 2397
rect 37921 2397 37933 2400
rect 37967 2397 37979 2431
rect 41417 2431 41475 2437
rect 41417 2428 41429 2431
rect 37921 2391 37979 2397
rect 38764 2400 41429 2428
rect 24762 2360 24768 2372
rect 23400 2332 24768 2360
rect 24762 2320 24768 2332
rect 24820 2320 24826 2372
rect 28353 2363 28411 2369
rect 28353 2329 28365 2363
rect 28399 2360 28411 2363
rect 30650 2360 30656 2372
rect 28399 2332 30656 2360
rect 28399 2329 28411 2332
rect 28353 2323 28411 2329
rect 30650 2320 30656 2332
rect 30708 2320 30714 2372
rect 37734 2320 37740 2372
rect 37792 2360 37798 2372
rect 38764 2360 38792 2400
rect 41417 2397 41429 2400
rect 41463 2397 41475 2431
rect 41417 2391 41475 2397
rect 42797 2431 42855 2437
rect 42797 2397 42809 2431
rect 42843 2397 42855 2431
rect 42797 2391 42855 2397
rect 37792 2332 38792 2360
rect 37792 2320 37798 2332
rect 40770 2320 40776 2372
rect 40828 2360 40834 2372
rect 42812 2360 42840 2391
rect 42978 2388 42984 2440
rect 43036 2428 43042 2440
rect 44821 2431 44879 2437
rect 44821 2428 44833 2431
rect 43036 2400 44833 2428
rect 43036 2388 43042 2400
rect 44821 2397 44833 2400
rect 44867 2397 44879 2431
rect 46201 2431 46259 2437
rect 46201 2428 46213 2431
rect 44821 2391 44879 2397
rect 45526 2400 46213 2428
rect 40828 2332 42840 2360
rect 40828 2320 40834 2332
rect 44358 2320 44364 2372
rect 44416 2360 44422 2372
rect 45526 2360 45554 2400
rect 46201 2397 46213 2400
rect 46247 2397 46259 2431
rect 46201 2391 46259 2397
rect 47581 2431 47639 2437
rect 47581 2397 47593 2431
rect 47627 2397 47639 2431
rect 47581 2391 47639 2397
rect 44416 2332 45554 2360
rect 44416 2320 44422 2332
rect 45738 2320 45744 2372
rect 45796 2360 45802 2372
rect 47596 2360 47624 2391
rect 48498 2388 48504 2440
rect 48556 2428 48562 2440
rect 50341 2431 50399 2437
rect 50341 2428 50353 2431
rect 48556 2400 50353 2428
rect 48556 2388 48562 2400
rect 50341 2397 50353 2400
rect 50387 2397 50399 2431
rect 50341 2391 50399 2397
rect 52457 2431 52515 2437
rect 52457 2397 52469 2431
rect 52503 2397 52515 2431
rect 52457 2391 52515 2397
rect 45796 2332 47624 2360
rect 45796 2320 45802 2332
rect 50706 2320 50712 2372
rect 50764 2360 50770 2372
rect 52472 2360 52500 2391
rect 50764 2332 52500 2360
rect 50764 2320 50770 2332
rect 22738 2252 22744 2304
rect 22796 2292 22802 2304
rect 25866 2292 25872 2304
rect 22796 2264 25872 2292
rect 22796 2252 22802 2264
rect 25866 2252 25872 2264
rect 25924 2252 25930 2304
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 19978 2048 19984 2100
rect 20036 2088 20042 2100
rect 23658 2088 23664 2100
rect 20036 2060 23664 2088
rect 20036 2048 20042 2060
rect 23658 2048 23664 2060
rect 23716 2048 23722 2100
rect 21358 1980 21364 2032
rect 21416 2020 21422 2032
rect 25314 2020 25320 2032
rect 21416 1992 25320 2020
rect 21416 1980 21422 1992
rect 25314 1980 25320 1992
rect 25372 1980 25378 2032
rect 24854 1368 24860 1420
rect 24912 1408 24918 1420
rect 25590 1408 25596 1420
rect 24912 1380 25596 1408
rect 24912 1368 24918 1380
rect 25590 1368 25596 1380
rect 25648 1368 25654 1420
<< via1 >>
rect 20168 57876 20220 57928
rect 25412 57876 25464 57928
rect 27712 57876 27764 57928
rect 34704 57876 34756 57928
rect 39120 57876 39172 57928
rect 43444 57876 43496 57928
rect 21824 57808 21876 57860
rect 26424 57808 26476 57860
rect 28080 57808 28132 57860
rect 36176 57808 36228 57860
rect 40132 57808 40184 57860
rect 51264 57808 51316 57860
rect 13268 57740 13320 57792
rect 24216 57740 24268 57792
rect 24492 57740 24544 57792
rect 39948 57740 40000 57792
rect 40500 57740 40552 57792
rect 44824 57740 44876 57792
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 3700 57536 3752 57588
rect 5540 57536 5592 57588
rect 10600 57536 10652 57588
rect 11980 57536 12032 57588
rect 13360 57536 13412 57588
rect 14740 57536 14792 57588
rect 16120 57536 16172 57588
rect 17500 57536 17552 57588
rect 18880 57536 18932 57588
rect 20260 57536 20312 57588
rect 21548 57536 21600 57588
rect 24400 57536 24452 57588
rect 29000 57536 29052 57588
rect 29644 57536 29696 57588
rect 30288 57536 30340 57588
rect 6368 57443 6420 57452
rect 6368 57409 6377 57443
rect 6377 57409 6411 57443
rect 6411 57409 6420 57443
rect 6368 57400 6420 57409
rect 7380 57400 7432 57452
rect 8300 57443 8352 57452
rect 8300 57409 8309 57443
rect 8309 57409 8343 57443
rect 8343 57409 8352 57443
rect 8300 57400 8352 57409
rect 9220 57400 9272 57452
rect 11888 57443 11940 57452
rect 11060 57264 11112 57316
rect 11888 57409 11897 57443
rect 11897 57409 11931 57443
rect 11931 57409 11940 57443
rect 11888 57400 11940 57409
rect 13268 57443 13320 57452
rect 13268 57409 13277 57443
rect 13277 57409 13311 57443
rect 13311 57409 13320 57443
rect 13268 57400 13320 57409
rect 21456 57468 21508 57520
rect 21732 57468 21784 57520
rect 26976 57468 27028 57520
rect 27160 57468 27212 57520
rect 17408 57443 17460 57452
rect 17408 57409 17417 57443
rect 17417 57409 17451 57443
rect 17451 57409 17460 57443
rect 17408 57400 17460 57409
rect 20168 57443 20220 57452
rect 20168 57409 20177 57443
rect 20177 57409 20211 57443
rect 20211 57409 20220 57443
rect 20168 57400 20220 57409
rect 21824 57400 21876 57452
rect 21916 57400 21968 57452
rect 22284 57332 22336 57384
rect 23756 57400 23808 57452
rect 24124 57443 24176 57452
rect 24124 57409 24133 57443
rect 24133 57409 24167 57443
rect 24167 57409 24176 57443
rect 24124 57400 24176 57409
rect 24308 57443 24360 57452
rect 24308 57409 24317 57443
rect 24317 57409 24351 57443
rect 24351 57409 24360 57443
rect 24308 57400 24360 57409
rect 25228 57400 25280 57452
rect 25504 57443 25556 57452
rect 25504 57409 25513 57443
rect 25513 57409 25547 57443
rect 25547 57409 25556 57443
rect 25504 57400 25556 57409
rect 23664 57332 23716 57384
rect 25044 57264 25096 57316
rect 20720 57196 20772 57248
rect 21916 57196 21968 57248
rect 22100 57239 22152 57248
rect 22100 57205 22109 57239
rect 22109 57205 22143 57239
rect 22143 57205 22152 57239
rect 26240 57332 26292 57384
rect 26884 57443 26936 57452
rect 26884 57409 26893 57443
rect 26893 57409 26927 57443
rect 26927 57409 26936 57443
rect 26884 57400 26936 57409
rect 27712 57400 27764 57452
rect 27896 57443 27948 57452
rect 27896 57409 27905 57443
rect 27905 57409 27939 57443
rect 27939 57409 27948 57443
rect 27896 57400 27948 57409
rect 28172 57468 28224 57520
rect 30656 57536 30708 57588
rect 35532 57536 35584 57588
rect 39948 57536 40000 57588
rect 43812 57536 43864 57588
rect 43996 57536 44048 57588
rect 51264 57579 51316 57588
rect 32956 57468 33008 57520
rect 27620 57375 27672 57384
rect 27620 57341 27629 57375
rect 27629 57341 27663 57375
rect 27663 57341 27672 57375
rect 27620 57332 27672 57341
rect 28172 57332 28224 57384
rect 29460 57400 29512 57452
rect 31760 57443 31812 57452
rect 31760 57409 31769 57443
rect 31769 57409 31803 57443
rect 31803 57409 31812 57443
rect 31760 57400 31812 57409
rect 33692 57400 33744 57452
rect 33784 57400 33836 57452
rect 35624 57468 35676 57520
rect 34796 57400 34848 57452
rect 36268 57400 36320 57452
rect 40224 57468 40276 57520
rect 38660 57443 38712 57452
rect 38660 57409 38669 57443
rect 38669 57409 38703 57443
rect 38703 57409 38712 57443
rect 38660 57400 38712 57409
rect 39856 57400 39908 57452
rect 45560 57468 45612 57520
rect 45836 57511 45888 57520
rect 45836 57477 45845 57511
rect 45845 57477 45879 57511
rect 45879 57477 45888 57511
rect 45836 57468 45888 57477
rect 46940 57443 46992 57452
rect 32404 57332 32456 57384
rect 35900 57375 35952 57384
rect 35900 57341 35909 57375
rect 35909 57341 35943 57375
rect 35943 57341 35952 57375
rect 35900 57332 35952 57341
rect 37280 57375 37332 57384
rect 37280 57341 37289 57375
rect 37289 57341 37323 57375
rect 37323 57341 37332 57375
rect 37280 57332 37332 57341
rect 37464 57332 37516 57384
rect 28264 57264 28316 57316
rect 28908 57264 28960 57316
rect 33416 57264 33468 57316
rect 22100 57196 22152 57205
rect 25596 57196 25648 57248
rect 27068 57239 27120 57248
rect 27068 57205 27077 57239
rect 27077 57205 27111 57239
rect 27111 57205 27120 57239
rect 27068 57196 27120 57205
rect 27712 57239 27764 57248
rect 27712 57205 27721 57239
rect 27721 57205 27755 57239
rect 27755 57205 27764 57239
rect 27712 57196 27764 57205
rect 29276 57196 29328 57248
rect 29368 57196 29420 57248
rect 30656 57196 30708 57248
rect 31024 57196 31076 57248
rect 32220 57196 32272 57248
rect 34336 57196 34388 57248
rect 34612 57264 34664 57316
rect 40316 57375 40368 57384
rect 40316 57341 40325 57375
rect 40325 57341 40359 57375
rect 40359 57341 40368 57375
rect 40316 57332 40368 57341
rect 40500 57375 40552 57384
rect 40500 57341 40509 57375
rect 40509 57341 40543 57375
rect 40543 57341 40552 57375
rect 40500 57332 40552 57341
rect 42892 57332 42944 57384
rect 43076 57375 43128 57384
rect 43076 57341 43085 57375
rect 43085 57341 43119 57375
rect 43119 57341 43128 57375
rect 43076 57332 43128 57341
rect 43812 57332 43864 57384
rect 46940 57409 46949 57443
rect 46949 57409 46983 57443
rect 46983 57409 46992 57443
rect 46940 57400 46992 57409
rect 48320 57443 48372 57452
rect 48320 57409 48329 57443
rect 48329 57409 48363 57443
rect 48363 57409 48372 57443
rect 48320 57400 48372 57409
rect 51264 57545 51273 57579
rect 51273 57545 51307 57579
rect 51307 57545 51316 57579
rect 51264 57536 51316 57545
rect 52460 57536 52512 57588
rect 52552 57468 52604 57520
rect 49700 57443 49752 57452
rect 49700 57409 49709 57443
rect 49709 57409 49743 57443
rect 49743 57409 49752 57443
rect 49700 57400 49752 57409
rect 51080 57400 51132 57452
rect 51632 57400 51684 57452
rect 53840 57400 53892 57452
rect 55220 57400 55272 57452
rect 55680 57400 55732 57452
rect 40592 57264 40644 57316
rect 36452 57196 36504 57248
rect 40132 57196 40184 57248
rect 40776 57196 40828 57248
rect 44180 57239 44232 57248
rect 44180 57205 44189 57239
rect 44189 57205 44223 57239
rect 44223 57205 44232 57239
rect 44180 57196 44232 57205
rect 44548 57332 44600 57384
rect 44732 57332 44784 57384
rect 47216 57375 47268 57384
rect 47216 57341 47225 57375
rect 47225 57341 47259 57375
rect 47259 57341 47268 57375
rect 47216 57332 47268 57341
rect 50068 57264 50120 57316
rect 45008 57196 45060 57248
rect 45744 57239 45796 57248
rect 45744 57205 45753 57239
rect 45753 57205 45787 57239
rect 45787 57205 45796 57239
rect 45744 57196 45796 57205
rect 51080 57196 51132 57248
rect 54116 57239 54168 57248
rect 54116 57205 54125 57239
rect 54125 57205 54159 57239
rect 54159 57205 54168 57239
rect 54116 57196 54168 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 4620 56992 4672 57044
rect 6000 56992 6052 57044
rect 6460 56992 6512 57044
rect 8760 56992 8812 57044
rect 10140 56992 10192 57044
rect 11520 56992 11572 57044
rect 12900 56992 12952 57044
rect 14280 56992 14332 57044
rect 15660 56992 15712 57044
rect 17040 56992 17092 57044
rect 18420 56992 18472 57044
rect 19984 56992 20036 57044
rect 21180 56992 21232 57044
rect 23020 57035 23072 57044
rect 23020 57001 23029 57035
rect 23029 57001 23063 57035
rect 23063 57001 23072 57035
rect 23020 56992 23072 57001
rect 24216 56992 24268 57044
rect 26976 56992 27028 57044
rect 28080 57035 28132 57044
rect 28080 57001 28089 57035
rect 28089 57001 28123 57035
rect 28123 57001 28132 57035
rect 28080 56992 28132 57001
rect 28172 56992 28224 57044
rect 32680 56992 32732 57044
rect 22284 56967 22336 56976
rect 22284 56933 22293 56967
rect 22293 56933 22327 56967
rect 22327 56933 22336 56967
rect 22284 56924 22336 56933
rect 27988 56924 28040 56976
rect 28448 56924 28500 56976
rect 28908 56924 28960 56976
rect 11060 56856 11112 56908
rect 22100 56856 22152 56908
rect 25412 56856 25464 56908
rect 23204 56831 23256 56840
rect 23204 56797 23213 56831
rect 23213 56797 23247 56831
rect 23247 56797 23256 56831
rect 23204 56788 23256 56797
rect 23756 56831 23808 56840
rect 23756 56797 23765 56831
rect 23765 56797 23799 56831
rect 23799 56797 23808 56831
rect 23756 56788 23808 56797
rect 24124 56788 24176 56840
rect 24032 56720 24084 56772
rect 25504 56788 25556 56840
rect 25872 56856 25924 56908
rect 26424 56899 26476 56908
rect 26424 56865 26433 56899
rect 26433 56865 26467 56899
rect 26467 56865 26476 56899
rect 26424 56856 26476 56865
rect 26516 56899 26568 56908
rect 26516 56865 26525 56899
rect 26525 56865 26559 56899
rect 26559 56865 26568 56899
rect 26516 56856 26568 56865
rect 27160 56856 27212 56908
rect 27712 56856 27764 56908
rect 27344 56788 27396 56840
rect 27436 56788 27488 56840
rect 27528 56720 27580 56772
rect 29184 56856 29236 56908
rect 29368 56924 29420 56976
rect 29552 56924 29604 56976
rect 37372 56992 37424 57044
rect 28172 56831 28224 56840
rect 28172 56797 28181 56831
rect 28181 56797 28215 56831
rect 28215 56797 28224 56831
rect 28172 56788 28224 56797
rect 29276 56831 29328 56840
rect 29276 56797 29285 56831
rect 29285 56797 29319 56831
rect 29319 56797 29328 56831
rect 29276 56788 29328 56797
rect 29368 56788 29420 56840
rect 29828 56831 29880 56840
rect 28080 56720 28132 56772
rect 28540 56720 28592 56772
rect 29828 56797 29837 56831
rect 29837 56797 29871 56831
rect 29871 56797 29880 56831
rect 29828 56788 29880 56797
rect 34796 56924 34848 56976
rect 31024 56831 31076 56840
rect 31024 56797 31033 56831
rect 31033 56797 31067 56831
rect 31067 56797 31076 56831
rect 31024 56788 31076 56797
rect 31760 56788 31812 56840
rect 33416 56831 33468 56840
rect 24492 56652 24544 56704
rect 25044 56652 25096 56704
rect 25504 56652 25556 56704
rect 26884 56695 26936 56704
rect 26884 56661 26893 56695
rect 26893 56661 26927 56695
rect 26927 56661 26936 56695
rect 26884 56652 26936 56661
rect 29460 56652 29512 56704
rect 30012 56652 30064 56704
rect 31760 56695 31812 56704
rect 31760 56661 31769 56695
rect 31769 56661 31803 56695
rect 31803 56661 31812 56695
rect 32220 56720 32272 56772
rect 33416 56797 33425 56831
rect 33425 56797 33459 56831
rect 33459 56797 33468 56831
rect 33416 56788 33468 56797
rect 34336 56856 34388 56908
rect 33784 56831 33836 56840
rect 33784 56797 33793 56831
rect 33793 56797 33827 56831
rect 33827 56797 33836 56831
rect 34428 56831 34480 56840
rect 33784 56788 33836 56797
rect 34428 56797 34437 56831
rect 34437 56797 34471 56831
rect 34471 56797 34480 56831
rect 34428 56788 34480 56797
rect 34612 56831 34664 56840
rect 34612 56797 34621 56831
rect 34621 56797 34655 56831
rect 34655 56797 34664 56831
rect 34612 56788 34664 56797
rect 34888 56788 34940 56840
rect 36452 56720 36504 56772
rect 31760 56652 31812 56661
rect 32036 56652 32088 56704
rect 33232 56695 33284 56704
rect 33232 56661 33241 56695
rect 33241 56661 33275 56695
rect 33275 56661 33284 56695
rect 33232 56652 33284 56661
rect 36084 56695 36136 56704
rect 36084 56661 36093 56695
rect 36093 56661 36127 56695
rect 36127 56661 36136 56695
rect 36084 56652 36136 56661
rect 37280 56788 37332 56840
rect 37832 56856 37884 56908
rect 39764 56924 39816 56976
rect 40408 56924 40460 56976
rect 43812 56924 43864 56976
rect 46020 56992 46072 57044
rect 48780 56992 48832 57044
rect 49700 57035 49752 57044
rect 49700 57001 49709 57035
rect 49709 57001 49743 57035
rect 49743 57001 49752 57035
rect 49700 56992 49752 57001
rect 50160 56992 50212 57044
rect 50620 56992 50672 57044
rect 51540 56992 51592 57044
rect 52460 57035 52512 57044
rect 52460 57001 52469 57035
rect 52469 57001 52503 57035
rect 52503 57001 52512 57035
rect 52460 56992 52512 57001
rect 52920 56992 52972 57044
rect 53380 56992 53432 57044
rect 54300 56992 54352 57044
rect 56140 56992 56192 57044
rect 46940 56924 46992 56976
rect 38844 56831 38896 56840
rect 38844 56797 38853 56831
rect 38853 56797 38887 56831
rect 38887 56797 38896 56831
rect 38844 56788 38896 56797
rect 38936 56831 38988 56840
rect 38936 56797 38945 56831
rect 38945 56797 38979 56831
rect 38979 56797 38988 56831
rect 38936 56788 38988 56797
rect 40132 56788 40184 56840
rect 40224 56788 40276 56840
rect 44180 56899 44232 56908
rect 41788 56831 41840 56840
rect 41788 56797 41797 56831
rect 41797 56797 41831 56831
rect 41831 56797 41840 56831
rect 41788 56788 41840 56797
rect 42708 56831 42760 56840
rect 42708 56797 42717 56831
rect 42717 56797 42751 56831
rect 42751 56797 42760 56831
rect 42708 56788 42760 56797
rect 43444 56831 43496 56840
rect 43444 56797 43453 56831
rect 43453 56797 43487 56831
rect 43487 56797 43496 56831
rect 43444 56788 43496 56797
rect 44180 56865 44189 56899
rect 44189 56865 44223 56899
rect 44223 56865 44232 56899
rect 44180 56856 44232 56865
rect 45008 56899 45060 56908
rect 45008 56865 45017 56899
rect 45017 56865 45051 56899
rect 45051 56865 45060 56899
rect 54116 56924 54168 56976
rect 45008 56856 45060 56865
rect 54760 56856 54812 56908
rect 44088 56788 44140 56840
rect 44732 56831 44784 56840
rect 42156 56720 42208 56772
rect 44732 56797 44741 56831
rect 44741 56797 44775 56831
rect 44775 56797 44784 56831
rect 44732 56788 44784 56797
rect 45652 56831 45704 56840
rect 45652 56797 45661 56831
rect 45661 56797 45695 56831
rect 45695 56797 45704 56831
rect 45652 56788 45704 56797
rect 46112 56831 46164 56840
rect 46112 56797 46121 56831
rect 46121 56797 46155 56831
rect 46155 56797 46164 56831
rect 46112 56788 46164 56797
rect 46940 56831 46992 56840
rect 46940 56797 46949 56831
rect 46949 56797 46983 56831
rect 46983 56797 46992 56831
rect 46940 56788 46992 56797
rect 40316 56652 40368 56704
rect 40592 56652 40644 56704
rect 41328 56652 41380 56704
rect 43168 56652 43220 56704
rect 45468 56695 45520 56704
rect 45468 56661 45477 56695
rect 45477 56661 45511 56695
rect 45511 56661 45520 56695
rect 45468 56652 45520 56661
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 24032 56491 24084 56500
rect 24032 56457 24041 56491
rect 24041 56457 24075 56491
rect 24075 56457 24084 56491
rect 24032 56448 24084 56457
rect 28172 56448 28224 56500
rect 27896 56380 27948 56432
rect 28632 56380 28684 56432
rect 22560 56312 22612 56364
rect 24492 56312 24544 56364
rect 25504 56355 25556 56364
rect 25504 56321 25513 56355
rect 25513 56321 25547 56355
rect 25547 56321 25556 56355
rect 25504 56312 25556 56321
rect 26240 56355 26292 56364
rect 26240 56321 26259 56355
rect 26259 56321 26292 56355
rect 27344 56355 27396 56364
rect 26240 56312 26292 56321
rect 27344 56321 27353 56355
rect 27353 56321 27387 56355
rect 27387 56321 27396 56355
rect 27344 56312 27396 56321
rect 28264 56355 28316 56364
rect 28264 56321 28273 56355
rect 28273 56321 28307 56355
rect 28307 56321 28316 56355
rect 28264 56312 28316 56321
rect 23664 56244 23716 56296
rect 25136 56244 25188 56296
rect 27712 56244 27764 56296
rect 27988 56244 28040 56296
rect 30472 56448 30524 56500
rect 31852 56448 31904 56500
rect 32680 56491 32732 56500
rect 32680 56457 32689 56491
rect 32689 56457 32723 56491
rect 32723 56457 32732 56491
rect 32680 56448 32732 56457
rect 30748 56380 30800 56432
rect 34520 56448 34572 56500
rect 34796 56448 34848 56500
rect 35532 56491 35584 56500
rect 35532 56457 35541 56491
rect 35541 56457 35575 56491
rect 35575 56457 35584 56491
rect 35532 56448 35584 56457
rect 36176 56448 36228 56500
rect 37280 56491 37332 56500
rect 37280 56457 37289 56491
rect 37289 56457 37323 56491
rect 37323 56457 37332 56491
rect 37280 56448 37332 56457
rect 29368 56355 29420 56364
rect 29368 56321 29377 56355
rect 29377 56321 29411 56355
rect 29411 56321 29420 56355
rect 29368 56312 29420 56321
rect 29460 56355 29512 56364
rect 29460 56321 29469 56355
rect 29469 56321 29503 56355
rect 29503 56321 29512 56355
rect 29460 56312 29512 56321
rect 23204 56176 23256 56228
rect 29276 56219 29328 56228
rect 29276 56185 29285 56219
rect 29285 56185 29319 56219
rect 29319 56185 29328 56219
rect 29276 56176 29328 56185
rect 29828 56312 29880 56364
rect 30196 56312 30248 56364
rect 30840 56312 30892 56364
rect 31760 56312 31812 56364
rect 32220 56355 32272 56364
rect 32220 56321 32229 56355
rect 32229 56321 32263 56355
rect 32263 56321 32272 56355
rect 32220 56312 32272 56321
rect 33232 56312 33284 56364
rect 30472 56287 30524 56296
rect 30472 56253 30481 56287
rect 30481 56253 30515 56287
rect 30515 56253 30524 56287
rect 30472 56244 30524 56253
rect 33140 56287 33192 56296
rect 33140 56253 33149 56287
rect 33149 56253 33183 56287
rect 33183 56253 33192 56287
rect 33140 56244 33192 56253
rect 33692 56176 33744 56228
rect 25688 56151 25740 56160
rect 25688 56117 25697 56151
rect 25697 56117 25731 56151
rect 25731 56117 25740 56151
rect 25688 56108 25740 56117
rect 27160 56151 27212 56160
rect 27160 56117 27169 56151
rect 27169 56117 27203 56151
rect 27203 56117 27212 56151
rect 27160 56108 27212 56117
rect 29000 56151 29052 56160
rect 29000 56117 29009 56151
rect 29009 56117 29043 56151
rect 29043 56117 29052 56151
rect 29000 56108 29052 56117
rect 30104 56151 30156 56160
rect 30104 56117 30113 56151
rect 30113 56117 30147 56151
rect 30147 56117 30156 56151
rect 30104 56108 30156 56117
rect 31852 56108 31904 56160
rect 32036 56108 32088 56160
rect 33048 56151 33100 56160
rect 33048 56117 33057 56151
rect 33057 56117 33091 56151
rect 33091 56117 33100 56151
rect 33048 56108 33100 56117
rect 34704 56423 34756 56432
rect 34704 56389 34713 56423
rect 34713 56389 34747 56423
rect 34747 56389 34756 56423
rect 34704 56380 34756 56389
rect 34888 56380 34940 56432
rect 34612 56312 34664 56364
rect 33876 56108 33928 56160
rect 33968 56108 34020 56160
rect 35532 56312 35584 56364
rect 37832 56380 37884 56432
rect 40776 56380 40828 56432
rect 37648 56355 37700 56364
rect 37648 56321 37657 56355
rect 37657 56321 37691 56355
rect 37691 56321 37700 56355
rect 37648 56312 37700 56321
rect 38844 56312 38896 56364
rect 39212 56355 39264 56364
rect 39212 56321 39221 56355
rect 39221 56321 39255 56355
rect 39255 56321 39264 56355
rect 39212 56312 39264 56321
rect 38568 56244 38620 56296
rect 36176 56108 36228 56160
rect 38108 56176 38160 56228
rect 38936 56176 38988 56228
rect 39764 56312 39816 56364
rect 40132 56312 40184 56364
rect 40040 56287 40092 56296
rect 40040 56253 40049 56287
rect 40049 56253 40083 56287
rect 40083 56253 40092 56287
rect 40040 56244 40092 56253
rect 40960 56312 41012 56364
rect 41328 56312 41380 56364
rect 42064 56448 42116 56500
rect 48320 56448 48372 56500
rect 49792 56448 49844 56500
rect 51632 56491 51684 56500
rect 51632 56457 51641 56491
rect 51641 56457 51675 56491
rect 51675 56457 51684 56491
rect 51632 56448 51684 56457
rect 52552 56448 52604 56500
rect 53840 56491 53892 56500
rect 53840 56457 53849 56491
rect 53849 56457 53883 56491
rect 53883 56457 53892 56491
rect 53840 56448 53892 56457
rect 55220 56491 55272 56500
rect 55220 56457 55229 56491
rect 55229 56457 55263 56491
rect 55263 56457 55272 56491
rect 55220 56448 55272 56457
rect 44088 56380 44140 56432
rect 45744 56380 45796 56432
rect 42156 56355 42208 56364
rect 42156 56321 42165 56355
rect 42165 56321 42199 56355
rect 42199 56321 42208 56355
rect 42156 56312 42208 56321
rect 43168 56355 43220 56364
rect 40408 56244 40460 56296
rect 40684 56219 40736 56228
rect 40684 56185 40693 56219
rect 40693 56185 40727 56219
rect 40727 56185 40736 56219
rect 40684 56176 40736 56185
rect 42800 56219 42852 56228
rect 42800 56185 42809 56219
rect 42809 56185 42843 56219
rect 42843 56185 42852 56219
rect 42800 56176 42852 56185
rect 43168 56321 43177 56355
rect 43177 56321 43211 56355
rect 43211 56321 43220 56355
rect 43168 56312 43220 56321
rect 43720 56312 43772 56364
rect 42984 56244 43036 56296
rect 43996 56355 44048 56364
rect 43996 56321 44005 56355
rect 44005 56321 44039 56355
rect 44039 56321 44048 56355
rect 43996 56312 44048 56321
rect 44364 56312 44416 56364
rect 44824 56355 44876 56364
rect 44824 56321 44833 56355
rect 44833 56321 44867 56355
rect 44867 56321 44876 56355
rect 44824 56312 44876 56321
rect 45100 56312 45152 56364
rect 47400 56312 47452 56364
rect 47860 56312 47912 56364
rect 45560 56287 45612 56296
rect 43720 56176 43772 56228
rect 44088 56219 44140 56228
rect 44088 56185 44097 56219
rect 44097 56185 44131 56219
rect 44131 56185 44140 56219
rect 44088 56176 44140 56185
rect 44180 56219 44232 56228
rect 44180 56185 44189 56219
rect 44189 56185 44223 56219
rect 44223 56185 44232 56219
rect 45560 56253 45569 56287
rect 45569 56253 45603 56287
rect 45603 56253 45612 56287
rect 45560 56244 45612 56253
rect 44180 56176 44232 56185
rect 41144 56151 41196 56160
rect 41144 56117 41153 56151
rect 41153 56117 41187 56151
rect 41187 56117 41196 56151
rect 41144 56108 41196 56117
rect 41604 56108 41656 56160
rect 42708 56108 42760 56160
rect 44824 56108 44876 56160
rect 47216 56108 47268 56160
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 23664 55947 23716 55956
rect 23664 55913 23673 55947
rect 23673 55913 23707 55947
rect 23707 55913 23716 55947
rect 23664 55904 23716 55913
rect 23756 55904 23808 55956
rect 25780 55904 25832 55956
rect 17408 55836 17460 55888
rect 29000 55904 29052 55956
rect 30196 55904 30248 55956
rect 34428 55904 34480 55956
rect 39212 55947 39264 55956
rect 28264 55836 28316 55888
rect 28632 55879 28684 55888
rect 28632 55845 28641 55879
rect 28641 55845 28675 55879
rect 28675 55845 28684 55879
rect 28632 55836 28684 55845
rect 24308 55743 24360 55752
rect 24308 55709 24317 55743
rect 24317 55709 24351 55743
rect 24351 55709 24360 55743
rect 24308 55700 24360 55709
rect 27160 55768 27212 55820
rect 27528 55768 27580 55820
rect 33968 55836 34020 55888
rect 34060 55836 34112 55888
rect 35992 55836 36044 55888
rect 29184 55768 29236 55820
rect 30380 55768 30432 55820
rect 31024 55768 31076 55820
rect 25872 55743 25924 55752
rect 25872 55709 25881 55743
rect 25881 55709 25915 55743
rect 25915 55709 25924 55743
rect 25872 55700 25924 55709
rect 28816 55743 28868 55752
rect 27528 55632 27580 55684
rect 28816 55709 28825 55743
rect 28825 55709 28859 55743
rect 28859 55709 28868 55743
rect 28816 55700 28868 55709
rect 28908 55743 28960 55752
rect 28908 55709 28917 55743
rect 28917 55709 28951 55743
rect 28951 55709 28960 55743
rect 29644 55743 29696 55752
rect 28908 55700 28960 55709
rect 29644 55709 29653 55743
rect 29653 55709 29687 55743
rect 29687 55709 29696 55743
rect 29644 55700 29696 55709
rect 30288 55700 30340 55752
rect 34612 55811 34664 55820
rect 34612 55777 34621 55811
rect 34621 55777 34655 55811
rect 34655 55777 34664 55811
rect 34612 55768 34664 55777
rect 32128 55743 32180 55752
rect 32128 55709 32137 55743
rect 32137 55709 32171 55743
rect 32171 55709 32180 55743
rect 32128 55700 32180 55709
rect 32404 55743 32456 55752
rect 32404 55709 32413 55743
rect 32413 55709 32447 55743
rect 32447 55709 32456 55743
rect 32404 55700 32456 55709
rect 27988 55675 28040 55684
rect 27988 55641 27997 55675
rect 27997 55641 28031 55675
rect 28031 55641 28040 55675
rect 27988 55632 28040 55641
rect 30196 55632 30248 55684
rect 30932 55632 30984 55684
rect 33416 55700 33468 55752
rect 34704 55700 34756 55752
rect 36084 55768 36136 55820
rect 38016 55836 38068 55888
rect 38292 55836 38344 55888
rect 39212 55913 39221 55947
rect 39221 55913 39255 55947
rect 39255 55913 39264 55947
rect 39212 55904 39264 55913
rect 40500 55947 40552 55956
rect 40500 55913 40509 55947
rect 40509 55913 40543 55947
rect 40543 55913 40552 55947
rect 40500 55904 40552 55913
rect 40960 55904 41012 55956
rect 44364 55947 44416 55956
rect 44364 55913 44373 55947
rect 44373 55913 44407 55947
rect 44407 55913 44416 55947
rect 44364 55904 44416 55913
rect 44640 55904 44692 55956
rect 45836 55904 45888 55956
rect 47032 55904 47084 55956
rect 38568 55768 38620 55820
rect 37004 55743 37056 55752
rect 26516 55564 26568 55616
rect 28264 55564 28316 55616
rect 28908 55564 28960 55616
rect 29828 55607 29880 55616
rect 29828 55573 29837 55607
rect 29837 55573 29871 55607
rect 29871 55573 29880 55607
rect 29828 55564 29880 55573
rect 30012 55564 30064 55616
rect 33140 55564 33192 55616
rect 37004 55709 37013 55743
rect 37013 55709 37047 55743
rect 37047 55709 37056 55743
rect 37004 55700 37056 55709
rect 37648 55743 37700 55752
rect 37648 55709 37657 55743
rect 37657 55709 37691 55743
rect 37691 55709 37700 55743
rect 37648 55700 37700 55709
rect 36452 55632 36504 55684
rect 38292 55700 38344 55752
rect 37924 55632 37976 55684
rect 38936 55743 38988 55752
rect 38936 55709 38945 55743
rect 38945 55709 38979 55743
rect 38979 55709 38988 55743
rect 38936 55700 38988 55709
rect 39488 55700 39540 55752
rect 40592 55836 40644 55888
rect 40224 55768 40276 55820
rect 40316 55743 40368 55752
rect 40316 55709 40325 55743
rect 40325 55709 40359 55743
rect 40359 55709 40368 55743
rect 40316 55700 40368 55709
rect 44916 55836 44968 55888
rect 45100 55836 45152 55888
rect 51080 55836 51132 55888
rect 41788 55768 41840 55820
rect 41604 55743 41656 55752
rect 41604 55709 41613 55743
rect 41613 55709 41647 55743
rect 41647 55709 41656 55743
rect 41604 55700 41656 55709
rect 42248 55700 42300 55752
rect 42524 55743 42576 55752
rect 42524 55709 42533 55743
rect 42533 55709 42567 55743
rect 42567 55709 42576 55743
rect 42524 55700 42576 55709
rect 43352 55768 43404 55820
rect 43628 55700 43680 55752
rect 43812 55700 43864 55752
rect 42616 55632 42668 55684
rect 43076 55632 43128 55684
rect 36176 55564 36228 55616
rect 38936 55564 38988 55616
rect 41420 55607 41472 55616
rect 41420 55573 41429 55607
rect 41429 55573 41463 55607
rect 41463 55573 41472 55607
rect 41420 55564 41472 55573
rect 41972 55564 42024 55616
rect 43628 55564 43680 55616
rect 43720 55564 43772 55616
rect 45560 55700 45612 55752
rect 50068 55768 50120 55820
rect 44824 55564 44876 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 25412 55360 25464 55412
rect 27344 55360 27396 55412
rect 30012 55360 30064 55412
rect 30104 55360 30156 55412
rect 30288 55403 30340 55412
rect 30288 55369 30290 55403
rect 30290 55369 30324 55403
rect 30324 55369 30340 55403
rect 30288 55360 30340 55369
rect 30932 55360 30984 55412
rect 34612 55360 34664 55412
rect 25688 55267 25740 55276
rect 25688 55233 25697 55267
rect 25697 55233 25731 55267
rect 25731 55233 25740 55267
rect 25688 55224 25740 55233
rect 26240 55224 26292 55276
rect 29184 55224 29236 55276
rect 23940 55156 23992 55208
rect 25320 55156 25372 55208
rect 27804 55156 27856 55208
rect 28816 55156 28868 55208
rect 29368 55267 29420 55276
rect 29368 55233 29377 55267
rect 29377 55233 29411 55267
rect 29411 55233 29420 55267
rect 30472 55292 30524 55344
rect 32128 55292 32180 55344
rect 35624 55360 35676 55412
rect 37924 55360 37976 55412
rect 41788 55360 41840 55412
rect 42524 55360 42576 55412
rect 29368 55224 29420 55233
rect 30012 55224 30064 55276
rect 30380 55267 30432 55276
rect 30380 55233 30389 55267
rect 30389 55233 30423 55267
rect 30423 55233 30432 55267
rect 30380 55224 30432 55233
rect 30288 55156 30340 55208
rect 32220 55224 32272 55276
rect 32772 55224 32824 55276
rect 33140 55224 33192 55276
rect 33600 55224 33652 55276
rect 35440 55292 35492 55344
rect 36176 55224 36228 55276
rect 36820 55224 36872 55276
rect 37280 55224 37332 55276
rect 27620 55088 27672 55140
rect 28264 55131 28316 55140
rect 28264 55097 28273 55131
rect 28273 55097 28307 55131
rect 28307 55097 28316 55131
rect 28264 55088 28316 55097
rect 36268 55156 36320 55208
rect 28724 55020 28776 55072
rect 31852 55020 31904 55072
rect 32312 55063 32364 55072
rect 32312 55029 32321 55063
rect 32321 55029 32355 55063
rect 32355 55029 32364 55063
rect 32312 55020 32364 55029
rect 32772 55063 32824 55072
rect 32772 55029 32781 55063
rect 32781 55029 32815 55063
rect 32815 55029 32824 55063
rect 32772 55020 32824 55029
rect 33416 55020 33468 55072
rect 33876 55020 33928 55072
rect 35992 55088 36044 55140
rect 38752 55292 38804 55344
rect 43076 55292 43128 55344
rect 38752 55156 38804 55208
rect 40224 55267 40276 55276
rect 40224 55233 40233 55267
rect 40233 55233 40267 55267
rect 40267 55233 40276 55267
rect 40224 55224 40276 55233
rect 42524 55224 42576 55276
rect 43904 55224 43956 55276
rect 44364 55360 44416 55412
rect 44732 55403 44784 55412
rect 44732 55369 44741 55403
rect 44741 55369 44775 55403
rect 44775 55369 44784 55403
rect 44732 55360 44784 55369
rect 45560 55403 45612 55412
rect 45560 55369 45569 55403
rect 45569 55369 45603 55403
rect 45603 55369 45612 55403
rect 45560 55360 45612 55369
rect 45652 55360 45704 55412
rect 44272 55292 44324 55344
rect 44180 55267 44232 55276
rect 44180 55233 44189 55267
rect 44189 55233 44223 55267
rect 44223 55233 44232 55267
rect 44180 55224 44232 55233
rect 39028 55088 39080 55140
rect 42616 55156 42668 55208
rect 44088 55156 44140 55208
rect 35716 55020 35768 55072
rect 39672 55020 39724 55072
rect 40592 55020 40644 55072
rect 40776 55020 40828 55072
rect 42248 55063 42300 55072
rect 42248 55029 42257 55063
rect 42257 55029 42291 55063
rect 42291 55029 42300 55063
rect 42248 55020 42300 55029
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 25136 54859 25188 54868
rect 25136 54825 25145 54859
rect 25145 54825 25179 54859
rect 25179 54825 25188 54859
rect 25136 54816 25188 54825
rect 25872 54816 25924 54868
rect 26240 54816 26292 54868
rect 26424 54816 26476 54868
rect 29276 54816 29328 54868
rect 29920 54816 29972 54868
rect 30472 54816 30524 54868
rect 31300 54816 31352 54868
rect 29460 54748 29512 54800
rect 25596 54655 25648 54664
rect 25596 54621 25605 54655
rect 25605 54621 25639 54655
rect 25639 54621 25648 54655
rect 25596 54612 25648 54621
rect 27068 54655 27120 54664
rect 27068 54621 27077 54655
rect 27077 54621 27111 54655
rect 27111 54621 27120 54655
rect 27068 54612 27120 54621
rect 28448 54680 28500 54732
rect 28724 54723 28776 54732
rect 28724 54689 28733 54723
rect 28733 54689 28767 54723
rect 28767 54689 28776 54723
rect 28724 54680 28776 54689
rect 30196 54680 30248 54732
rect 33048 54748 33100 54800
rect 32312 54723 32364 54732
rect 32312 54689 32321 54723
rect 32321 54689 32355 54723
rect 32355 54689 32364 54723
rect 32312 54680 32364 54689
rect 33876 54723 33928 54732
rect 33876 54689 33885 54723
rect 33885 54689 33919 54723
rect 33919 54689 33928 54723
rect 33876 54680 33928 54689
rect 34888 54748 34940 54800
rect 36268 54816 36320 54868
rect 36360 54816 36412 54868
rect 38108 54859 38160 54868
rect 38108 54825 38117 54859
rect 38117 54825 38151 54859
rect 38151 54825 38160 54859
rect 38108 54816 38160 54825
rect 38936 54816 38988 54868
rect 40132 54816 40184 54868
rect 42064 54816 42116 54868
rect 43260 54816 43312 54868
rect 44272 54816 44324 54868
rect 39764 54748 39816 54800
rect 40316 54723 40368 54732
rect 40316 54689 40325 54723
rect 40325 54689 40359 54723
rect 40359 54689 40368 54723
rect 40316 54680 40368 54689
rect 28540 54612 28592 54664
rect 29000 54612 29052 54664
rect 30380 54544 30432 54596
rect 32772 54612 32824 54664
rect 32404 54544 32456 54596
rect 35624 54612 35676 54664
rect 35716 54612 35768 54664
rect 36176 54655 36228 54664
rect 36176 54621 36185 54655
rect 36185 54621 36219 54655
rect 36219 54621 36228 54655
rect 36176 54612 36228 54621
rect 37832 54612 37884 54664
rect 38016 54612 38068 54664
rect 38752 54612 38804 54664
rect 39028 54655 39080 54664
rect 39028 54621 39037 54655
rect 39037 54621 39071 54655
rect 39071 54621 39080 54655
rect 39028 54612 39080 54621
rect 39488 54655 39540 54664
rect 39488 54621 39497 54655
rect 39497 54621 39531 54655
rect 39531 54621 39540 54655
rect 39488 54612 39540 54621
rect 39672 54655 39724 54664
rect 39672 54621 39681 54655
rect 39681 54621 39715 54655
rect 39715 54621 39724 54655
rect 39672 54612 39724 54621
rect 40500 54655 40552 54664
rect 40500 54621 40509 54655
rect 40509 54621 40543 54655
rect 40543 54621 40552 54655
rect 40500 54612 40552 54621
rect 40776 54655 40828 54664
rect 40776 54621 40785 54655
rect 40785 54621 40819 54655
rect 40819 54621 40828 54655
rect 40776 54612 40828 54621
rect 41328 54612 41380 54664
rect 42524 54612 42576 54664
rect 42984 54655 43036 54664
rect 42984 54621 42993 54655
rect 42993 54621 43027 54655
rect 43027 54621 43036 54655
rect 42984 54612 43036 54621
rect 41420 54544 41472 54596
rect 43168 54544 43220 54596
rect 33324 54476 33376 54528
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 26240 54315 26292 54324
rect 26240 54281 26249 54315
rect 26249 54281 26283 54315
rect 26283 54281 26292 54315
rect 26240 54272 26292 54281
rect 29368 54272 29420 54324
rect 30012 54315 30064 54324
rect 30012 54281 30021 54315
rect 30021 54281 30055 54315
rect 30055 54281 30064 54315
rect 30012 54272 30064 54281
rect 30288 54272 30340 54324
rect 33140 54272 33192 54324
rect 33692 54272 33744 54324
rect 36452 54272 36504 54324
rect 39672 54272 39724 54324
rect 41328 54315 41380 54324
rect 41328 54281 41337 54315
rect 41337 54281 41371 54315
rect 41371 54281 41380 54315
rect 41328 54272 41380 54281
rect 42248 54272 42300 54324
rect 42892 54272 42944 54324
rect 29460 54204 29512 54256
rect 26700 54136 26752 54188
rect 28908 54136 28960 54188
rect 30196 54179 30248 54188
rect 30196 54145 30205 54179
rect 30205 54145 30239 54179
rect 30239 54145 30248 54179
rect 30196 54136 30248 54145
rect 30380 54179 30432 54188
rect 30380 54145 30389 54179
rect 30389 54145 30423 54179
rect 30423 54145 30432 54179
rect 30380 54136 30432 54145
rect 30748 54204 30800 54256
rect 33232 54247 33284 54256
rect 33232 54213 33241 54247
rect 33241 54213 33275 54247
rect 33275 54213 33284 54247
rect 33232 54204 33284 54213
rect 31024 54179 31076 54188
rect 31024 54145 31033 54179
rect 31033 54145 31067 54179
rect 31067 54145 31076 54179
rect 31024 54136 31076 54145
rect 32404 54179 32456 54188
rect 32404 54145 32413 54179
rect 32413 54145 32447 54179
rect 32447 54145 32456 54179
rect 32404 54136 32456 54145
rect 32956 54136 33008 54188
rect 33140 54136 33192 54188
rect 33324 54179 33376 54188
rect 33324 54145 33333 54179
rect 33333 54145 33367 54179
rect 33367 54145 33376 54179
rect 33324 54136 33376 54145
rect 33508 54136 33560 54188
rect 33968 54179 34020 54188
rect 33968 54145 33977 54179
rect 33977 54145 34011 54179
rect 34011 54145 34020 54179
rect 33968 54136 34020 54145
rect 36176 54204 36228 54256
rect 40408 54204 40460 54256
rect 41604 54204 41656 54256
rect 33416 54068 33468 54120
rect 34888 54179 34940 54188
rect 34888 54145 34897 54179
rect 34897 54145 34931 54179
rect 34931 54145 34940 54179
rect 34888 54136 34940 54145
rect 35348 54136 35400 54188
rect 37280 54179 37332 54188
rect 37280 54145 37289 54179
rect 37289 54145 37323 54179
rect 37323 54145 37332 54179
rect 37280 54136 37332 54145
rect 37740 54136 37792 54188
rect 38200 54136 38252 54188
rect 39580 54136 39632 54188
rect 40316 54179 40368 54188
rect 40316 54145 40325 54179
rect 40325 54145 40359 54179
rect 40359 54145 40368 54179
rect 40316 54136 40368 54145
rect 41420 54136 41472 54188
rect 43720 54136 43772 54188
rect 35716 54068 35768 54120
rect 31852 54000 31904 54052
rect 40040 54043 40092 54052
rect 40040 54009 40049 54043
rect 40049 54009 40083 54043
rect 40083 54009 40092 54043
rect 40040 54000 40092 54009
rect 27712 53975 27764 53984
rect 27712 53941 27721 53975
rect 27721 53941 27755 53975
rect 27755 53941 27764 53975
rect 27712 53932 27764 53941
rect 40500 53932 40552 53984
rect 41972 53975 42024 53984
rect 41972 53941 41981 53975
rect 41981 53941 42015 53975
rect 42015 53941 42024 53975
rect 41972 53932 42024 53941
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 28080 53771 28132 53780
rect 28080 53737 28089 53771
rect 28089 53737 28123 53771
rect 28123 53737 28132 53771
rect 28080 53728 28132 53737
rect 28908 53728 28960 53780
rect 29000 53728 29052 53780
rect 29736 53728 29788 53780
rect 31024 53728 31076 53780
rect 31944 53771 31996 53780
rect 31944 53737 31953 53771
rect 31953 53737 31987 53771
rect 31987 53737 31996 53771
rect 31944 53728 31996 53737
rect 33232 53728 33284 53780
rect 33968 53771 34020 53780
rect 33968 53737 33977 53771
rect 33977 53737 34011 53771
rect 34011 53737 34020 53771
rect 33968 53728 34020 53737
rect 34796 53728 34848 53780
rect 36084 53728 36136 53780
rect 37464 53728 37516 53780
rect 40408 53771 40460 53780
rect 40408 53737 40417 53771
rect 40417 53737 40451 53771
rect 40451 53737 40460 53771
rect 40408 53728 40460 53737
rect 33416 53660 33468 53712
rect 35900 53660 35952 53712
rect 39856 53703 39908 53712
rect 39856 53669 39865 53703
rect 39865 53669 39899 53703
rect 39899 53669 39908 53703
rect 39856 53660 39908 53669
rect 32588 53635 32640 53644
rect 32588 53601 32597 53635
rect 32597 53601 32631 53635
rect 32631 53601 32640 53635
rect 32588 53592 32640 53601
rect 35992 53592 36044 53644
rect 36452 53635 36504 53644
rect 36452 53601 36461 53635
rect 36461 53601 36495 53635
rect 36495 53601 36504 53635
rect 36452 53592 36504 53601
rect 29184 53524 29236 53576
rect 30012 53524 30064 53576
rect 33140 53524 33192 53576
rect 33324 53499 33376 53508
rect 33324 53465 33351 53499
rect 33351 53465 33376 53499
rect 33324 53456 33376 53465
rect 29368 53388 29420 53440
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 31024 53184 31076 53236
rect 32588 53227 32640 53236
rect 32588 53193 32597 53227
rect 32597 53193 32631 53227
rect 32631 53193 32640 53227
rect 32588 53184 32640 53193
rect 36084 53184 36136 53236
rect 40408 53184 40460 53236
rect 35532 53116 35584 53168
rect 34796 52980 34848 53032
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 35992 52640 36044 52692
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 27712 8032 27764 8084
rect 30840 8032 30892 8084
rect 29644 7828 29696 7880
rect 29552 7692 29604 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 26240 7352 26292 7404
rect 29644 7395 29696 7404
rect 29644 7361 29653 7395
rect 29653 7361 29687 7395
rect 29687 7361 29696 7395
rect 29644 7352 29696 7361
rect 32036 7395 32088 7404
rect 32036 7361 32045 7395
rect 32045 7361 32079 7395
rect 32079 7361 32088 7395
rect 32036 7352 32088 7361
rect 32956 7352 33008 7404
rect 27436 7191 27488 7200
rect 27436 7157 27445 7191
rect 27445 7157 27479 7191
rect 27479 7157 27488 7191
rect 27436 7148 27488 7157
rect 27988 7191 28040 7200
rect 27988 7157 27997 7191
rect 27997 7157 28031 7191
rect 28031 7157 28040 7191
rect 27988 7148 28040 7157
rect 29460 7148 29512 7200
rect 30196 7191 30248 7200
rect 30196 7157 30205 7191
rect 30205 7157 30239 7191
rect 30239 7157 30248 7191
rect 30196 7148 30248 7157
rect 30932 7148 30984 7200
rect 32312 7148 32364 7200
rect 33232 7148 33284 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 32036 6808 32088 6860
rect 25228 6740 25280 6792
rect 26240 6783 26292 6792
rect 26240 6749 26249 6783
rect 26249 6749 26283 6783
rect 26283 6749 26292 6783
rect 26240 6740 26292 6749
rect 26608 6740 26660 6792
rect 27620 6783 27672 6792
rect 27620 6749 27629 6783
rect 27629 6749 27663 6783
rect 27663 6749 27672 6783
rect 27620 6740 27672 6749
rect 29000 6740 29052 6792
rect 29276 6740 29328 6792
rect 29368 6740 29420 6792
rect 30840 6783 30892 6792
rect 30840 6749 30849 6783
rect 30849 6749 30883 6783
rect 30883 6749 30892 6783
rect 30840 6740 30892 6749
rect 31760 6783 31812 6792
rect 31760 6749 31769 6783
rect 31769 6749 31803 6783
rect 31803 6749 31812 6783
rect 31760 6740 31812 6749
rect 33140 6783 33192 6792
rect 29644 6672 29696 6724
rect 32036 6672 32088 6724
rect 33140 6749 33149 6783
rect 33149 6749 33183 6783
rect 33183 6749 33192 6783
rect 33140 6740 33192 6749
rect 33968 6783 34020 6792
rect 33968 6749 33977 6783
rect 33977 6749 34011 6783
rect 34011 6749 34020 6783
rect 33968 6740 34020 6749
rect 25136 6647 25188 6656
rect 25136 6613 25145 6647
rect 25145 6613 25179 6647
rect 25179 6613 25188 6647
rect 25136 6604 25188 6613
rect 26792 6604 26844 6656
rect 33416 6604 33468 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 25136 6400 25188 6452
rect 27712 6400 27764 6452
rect 26792 6375 26844 6384
rect 26792 6341 26801 6375
rect 26801 6341 26835 6375
rect 26835 6341 26844 6375
rect 26792 6332 26844 6341
rect 29460 6375 29512 6384
rect 29460 6341 29469 6375
rect 29469 6341 29503 6375
rect 29503 6341 29512 6375
rect 29460 6332 29512 6341
rect 32036 6375 32088 6384
rect 32036 6341 32045 6375
rect 32045 6341 32079 6375
rect 32079 6341 32088 6375
rect 32036 6332 32088 6341
rect 25688 6307 25740 6316
rect 25688 6273 25697 6307
rect 25697 6273 25731 6307
rect 25731 6273 25740 6307
rect 25688 6264 25740 6273
rect 29276 6307 29328 6316
rect 29276 6273 29285 6307
rect 29285 6273 29319 6307
rect 29319 6273 29328 6307
rect 29276 6264 29328 6273
rect 30840 6264 30892 6316
rect 32956 6264 33008 6316
rect 24860 6196 24912 6248
rect 27528 6239 27580 6248
rect 27528 6205 27537 6239
rect 27537 6205 27571 6239
rect 27571 6205 27580 6239
rect 27528 6196 27580 6205
rect 30012 6239 30064 6248
rect 30012 6205 30021 6239
rect 30021 6205 30055 6239
rect 30055 6205 30064 6239
rect 30012 6196 30064 6205
rect 33600 6128 33652 6180
rect 25412 6060 25464 6112
rect 32128 6060 32180 6112
rect 34796 6060 34848 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 26700 5763 26752 5772
rect 26700 5729 26709 5763
rect 26709 5729 26743 5763
rect 26743 5729 26752 5763
rect 26700 5720 26752 5729
rect 28632 5763 28684 5772
rect 28632 5729 28641 5763
rect 28641 5729 28675 5763
rect 28675 5729 28684 5763
rect 28632 5720 28684 5729
rect 31760 5788 31812 5840
rect 33968 5788 34020 5840
rect 30932 5763 30984 5772
rect 30932 5729 30941 5763
rect 30941 5729 30975 5763
rect 30975 5729 30984 5763
rect 30932 5720 30984 5729
rect 31668 5763 31720 5772
rect 31668 5729 31677 5763
rect 31677 5729 31711 5763
rect 31711 5729 31720 5763
rect 31668 5720 31720 5729
rect 33324 5763 33376 5772
rect 33324 5729 33333 5763
rect 33333 5729 33367 5763
rect 33367 5729 33376 5763
rect 33324 5720 33376 5729
rect 34796 5763 34848 5772
rect 34796 5729 34805 5763
rect 34805 5729 34839 5763
rect 34839 5729 34848 5763
rect 34796 5720 34848 5729
rect 23388 5652 23440 5704
rect 24308 5695 24360 5704
rect 24308 5661 24317 5695
rect 24317 5661 24351 5695
rect 24351 5661 24360 5695
rect 24308 5652 24360 5661
rect 24952 5652 25004 5704
rect 27896 5695 27948 5704
rect 27896 5661 27905 5695
rect 27905 5661 27939 5695
rect 27939 5661 27948 5695
rect 27896 5652 27948 5661
rect 25504 5584 25556 5636
rect 28080 5627 28132 5636
rect 28080 5593 28089 5627
rect 28089 5593 28123 5627
rect 28123 5593 28132 5627
rect 28080 5584 28132 5593
rect 24032 5516 24084 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 24308 5176 24360 5228
rect 26148 5244 26200 5296
rect 27436 5244 27488 5296
rect 30196 5244 30248 5296
rect 33416 5287 33468 5296
rect 33416 5253 33425 5287
rect 33425 5253 33459 5287
rect 33459 5253 33468 5287
rect 33416 5244 33468 5253
rect 37924 5244 37976 5296
rect 25688 5219 25740 5228
rect 25688 5185 25697 5219
rect 25697 5185 25731 5219
rect 25731 5185 25740 5219
rect 25688 5176 25740 5185
rect 26608 5219 26660 5228
rect 26608 5185 26617 5219
rect 26617 5185 26651 5219
rect 26651 5185 26660 5219
rect 26608 5176 26660 5185
rect 29368 5219 29420 5228
rect 29368 5185 29377 5219
rect 29377 5185 29411 5219
rect 29411 5185 29420 5219
rect 29368 5176 29420 5185
rect 33600 5219 33652 5228
rect 33600 5185 33609 5219
rect 33609 5185 33643 5219
rect 33643 5185 33652 5219
rect 33600 5176 33652 5185
rect 24860 5108 24912 5160
rect 27712 5151 27764 5160
rect 27712 5117 27721 5151
rect 27721 5117 27755 5151
rect 27755 5117 27764 5151
rect 27712 5108 27764 5117
rect 30380 5151 30432 5160
rect 30380 5117 30389 5151
rect 30389 5117 30423 5151
rect 30423 5117 30432 5151
rect 30380 5108 30432 5117
rect 31760 5151 31812 5160
rect 31760 5117 31769 5151
rect 31769 5117 31803 5151
rect 31803 5117 31812 5151
rect 34520 5151 34572 5160
rect 31760 5108 31812 5117
rect 34520 5117 34529 5151
rect 34529 5117 34563 5151
rect 34563 5117 34572 5151
rect 34520 5108 34572 5117
rect 37188 5108 37240 5160
rect 22560 4972 22612 5024
rect 27804 4972 27856 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 37188 4811 37240 4820
rect 37188 4777 37197 4811
rect 37197 4777 37231 4811
rect 37231 4777 37240 4811
rect 37188 4768 37240 4777
rect 23940 4700 23992 4752
rect 33232 4700 33284 4752
rect 25044 4632 25096 4684
rect 25228 4675 25280 4684
rect 25228 4641 25237 4675
rect 25237 4641 25271 4675
rect 25271 4641 25280 4675
rect 25228 4632 25280 4641
rect 25412 4675 25464 4684
rect 25412 4641 25421 4675
rect 25421 4641 25455 4675
rect 25455 4641 25464 4675
rect 25412 4632 25464 4641
rect 26240 4675 26292 4684
rect 26240 4641 26249 4675
rect 26249 4641 26283 4675
rect 26283 4641 26292 4675
rect 26240 4632 26292 4641
rect 27620 4675 27672 4684
rect 27620 4641 27629 4675
rect 27629 4641 27663 4675
rect 27663 4641 27672 4675
rect 27620 4632 27672 4641
rect 27804 4675 27856 4684
rect 27804 4641 27813 4675
rect 27813 4641 27847 4675
rect 27847 4641 27856 4675
rect 27804 4632 27856 4641
rect 28172 4675 28224 4684
rect 28172 4641 28181 4675
rect 28181 4641 28215 4675
rect 28215 4641 28224 4675
rect 28172 4632 28224 4641
rect 30748 4632 30800 4684
rect 33140 4675 33192 4684
rect 33140 4641 33149 4675
rect 33149 4641 33183 4675
rect 33183 4641 33192 4675
rect 33140 4632 33192 4641
rect 33600 4675 33652 4684
rect 33600 4641 33609 4675
rect 33609 4641 33643 4675
rect 33643 4641 33652 4675
rect 33600 4632 33652 4641
rect 20720 4607 20772 4616
rect 20720 4573 20729 4607
rect 20729 4573 20763 4607
rect 20763 4573 20772 4607
rect 20720 4564 20772 4573
rect 22008 4564 22060 4616
rect 23480 4564 23532 4616
rect 24308 4564 24360 4616
rect 30380 4607 30432 4616
rect 30380 4573 30389 4607
rect 30389 4573 30423 4607
rect 30423 4573 30432 4607
rect 30380 4564 30432 4573
rect 36360 4564 36412 4616
rect 36728 4607 36780 4616
rect 36728 4573 36737 4607
rect 36737 4573 36771 4607
rect 36771 4573 36780 4607
rect 36728 4564 36780 4573
rect 37832 4607 37884 4616
rect 37832 4573 37841 4607
rect 37841 4573 37875 4607
rect 37875 4573 37884 4607
rect 37832 4564 37884 4573
rect 30656 4496 30708 4548
rect 22652 4428 22704 4480
rect 26148 4428 26200 4480
rect 36176 4428 36228 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 36176 4199 36228 4208
rect 36176 4165 36185 4199
rect 36185 4165 36219 4199
rect 36219 4165 36228 4199
rect 36176 4156 36228 4165
rect 23480 4088 23532 4140
rect 25320 4088 25372 4140
rect 29000 4088 29052 4140
rect 32128 4131 32180 4140
rect 32128 4097 32137 4131
rect 32137 4097 32171 4131
rect 32171 4097 32180 4131
rect 32128 4088 32180 4097
rect 36360 4131 36412 4140
rect 36360 4097 36369 4131
rect 36369 4097 36403 4131
rect 36403 4097 36412 4131
rect 36360 4088 36412 4097
rect 22284 4020 22336 4072
rect 23848 4063 23900 4072
rect 23848 4029 23857 4063
rect 23857 4029 23891 4063
rect 23891 4029 23900 4063
rect 23848 4020 23900 4029
rect 22100 3952 22152 4004
rect 22192 3952 22244 4004
rect 17132 3884 17184 3936
rect 18420 3884 18472 3936
rect 20076 3884 20128 3936
rect 20352 3884 20404 3936
rect 22468 3884 22520 3936
rect 25136 3884 25188 3936
rect 26516 3952 26568 4004
rect 29552 4020 29604 4072
rect 29736 4063 29788 4072
rect 29736 4029 29745 4063
rect 29745 4029 29779 4063
rect 29779 4029 29788 4063
rect 29736 4020 29788 4029
rect 32312 4063 32364 4072
rect 32312 4029 32321 4063
rect 32321 4029 32355 4063
rect 32355 4029 32364 4063
rect 32312 4020 32364 4029
rect 32772 4063 32824 4072
rect 32772 4029 32781 4063
rect 32781 4029 32815 4063
rect 32815 4029 32824 4063
rect 32772 4020 32824 4029
rect 34060 4020 34112 4072
rect 35808 4020 35860 4072
rect 39120 4020 39172 4072
rect 29184 3952 29236 4004
rect 37556 3952 37608 4004
rect 39948 3952 40000 4004
rect 26976 3884 27028 3936
rect 37280 3927 37332 3936
rect 37280 3893 37289 3927
rect 37289 3893 37323 3927
rect 37323 3893 37332 3927
rect 37280 3884 37332 3893
rect 38292 3884 38344 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 22100 3680 22152 3732
rect 24952 3680 25004 3732
rect 25136 3680 25188 3732
rect 28080 3680 28132 3732
rect 36912 3680 36964 3732
rect 37832 3680 37884 3732
rect 21732 3612 21784 3664
rect 26148 3612 26200 3664
rect 21180 3544 21232 3596
rect 22468 3587 22520 3596
rect 22468 3553 22477 3587
rect 22477 3553 22511 3587
rect 22511 3553 22520 3587
rect 22468 3544 22520 3553
rect 22652 3587 22704 3596
rect 22652 3553 22661 3587
rect 22661 3553 22695 3587
rect 22695 3553 22704 3587
rect 22652 3544 22704 3553
rect 25044 3544 25096 3596
rect 27988 3587 28040 3596
rect 27988 3553 27997 3587
rect 27997 3553 28031 3587
rect 28031 3553 28040 3587
rect 27988 3544 28040 3553
rect 36176 3612 36228 3664
rect 40500 3612 40552 3664
rect 42708 3612 42760 3664
rect 28356 3544 28408 3596
rect 30840 3544 30892 3596
rect 32220 3544 32272 3596
rect 33692 3544 33744 3596
rect 38568 3544 38620 3596
rect 41328 3544 41380 3596
rect 10232 3476 10284 3528
rect 12164 3476 12216 3528
rect 12992 3476 13044 3528
rect 14096 3476 14148 3528
rect 14924 3476 14976 3528
rect 15752 3476 15804 3528
rect 16580 3476 16632 3528
rect 17868 3476 17920 3528
rect 18696 3476 18748 3528
rect 19248 3476 19300 3528
rect 22376 3476 22428 3528
rect 30564 3519 30616 3528
rect 30564 3485 30573 3519
rect 30573 3485 30607 3519
rect 30607 3485 30616 3519
rect 30564 3476 30616 3485
rect 33140 3519 33192 3528
rect 33140 3485 33149 3519
rect 33149 3485 33183 3519
rect 33183 3485 33192 3519
rect 33140 3476 33192 3485
rect 35900 3519 35952 3528
rect 35900 3485 35909 3519
rect 35909 3485 35943 3519
rect 35943 3485 35952 3519
rect 35900 3476 35952 3485
rect 24216 3408 24268 3460
rect 25412 3451 25464 3460
rect 22100 3340 22152 3392
rect 23480 3340 23532 3392
rect 25412 3417 25421 3451
rect 25421 3417 25455 3451
rect 25455 3417 25464 3451
rect 25412 3408 25464 3417
rect 28908 3408 28960 3460
rect 30380 3408 30432 3460
rect 33876 3408 33928 3460
rect 36084 3451 36136 3460
rect 36084 3417 36093 3451
rect 36093 3417 36127 3451
rect 36127 3417 36136 3451
rect 36084 3408 36136 3417
rect 36636 3408 36688 3460
rect 38844 3408 38896 3460
rect 41880 3408 41932 3460
rect 43536 3476 43588 3528
rect 44916 3476 44968 3528
rect 46296 3476 46348 3528
rect 47676 3476 47728 3528
rect 49056 3476 49108 3528
rect 50620 3476 50672 3528
rect 51816 3476 51868 3528
rect 26424 3340 26476 3392
rect 35532 3340 35584 3392
rect 40040 3340 40092 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 22192 3179 22244 3188
rect 22192 3145 22201 3179
rect 22201 3145 22235 3179
rect 22235 3145 22244 3179
rect 22192 3136 22244 3145
rect 24492 3136 24544 3188
rect 33048 3136 33100 3188
rect 33600 3136 33652 3188
rect 35348 3136 35400 3188
rect 39304 3136 39356 3188
rect 24032 3111 24084 3120
rect 18972 2932 19024 2984
rect 24032 3077 24041 3111
rect 24041 3077 24075 3111
rect 24075 3077 24084 3111
rect 24032 3068 24084 3077
rect 27252 3068 27304 3120
rect 34152 3068 34204 3120
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22100 3000 22152 3009
rect 22376 3000 22428 3052
rect 25044 2932 25096 2984
rect 26608 2975 26660 2984
rect 26608 2941 26617 2975
rect 26617 2941 26651 2975
rect 26651 2941 26660 2975
rect 26608 2932 26660 2941
rect 26792 2975 26844 2984
rect 26792 2941 26801 2975
rect 26801 2941 26835 2975
rect 26835 2941 26844 2975
rect 26792 2932 26844 2941
rect 19432 2864 19484 2916
rect 22744 2864 22796 2916
rect 8576 2796 8628 2848
rect 9312 2796 9364 2848
rect 9956 2839 10008 2848
rect 9956 2805 9965 2839
rect 9965 2805 9999 2839
rect 9999 2805 10008 2839
rect 9956 2796 10008 2805
rect 10784 2796 10836 2848
rect 11336 2796 11388 2848
rect 11612 2796 11664 2848
rect 12716 2839 12768 2848
rect 12716 2805 12725 2839
rect 12725 2805 12759 2839
rect 12759 2805 12768 2839
rect 12716 2796 12768 2805
rect 13544 2796 13596 2848
rect 14372 2796 14424 2848
rect 15200 2796 15252 2848
rect 16028 2796 16080 2848
rect 16304 2796 16356 2848
rect 17316 2796 17368 2848
rect 20904 2796 20956 2848
rect 25504 2864 25556 2916
rect 28540 2932 28592 2984
rect 29552 2975 29604 2984
rect 29552 2941 29561 2975
rect 29561 2941 29595 2975
rect 29595 2941 29604 2975
rect 29552 2932 29604 2941
rect 31116 2975 31168 2984
rect 31116 2941 31125 2975
rect 31125 2941 31159 2975
rect 31159 2941 31168 2975
rect 31116 2932 31168 2941
rect 31944 2975 31996 2984
rect 31944 2941 31953 2975
rect 31953 2941 31987 2975
rect 31987 2941 31996 2975
rect 31944 2932 31996 2941
rect 33416 2975 33468 2984
rect 33416 2941 33425 2975
rect 33425 2941 33459 2975
rect 33459 2941 33468 2975
rect 33416 2932 33468 2941
rect 33600 2975 33652 2984
rect 33600 2941 33609 2975
rect 33609 2941 33643 2975
rect 33643 2941 33652 2975
rect 33600 2932 33652 2941
rect 34520 2975 34572 2984
rect 34520 2941 34529 2975
rect 34529 2941 34563 2975
rect 34563 2941 34572 2975
rect 34520 2932 34572 2941
rect 34704 2975 34756 2984
rect 34704 2941 34713 2975
rect 34713 2941 34747 2975
rect 34747 2941 34756 2975
rect 34704 2932 34756 2941
rect 29460 2864 29512 2916
rect 32496 2864 32548 2916
rect 36360 3068 36412 3120
rect 37280 3043 37332 3052
rect 37280 3009 37289 3043
rect 37289 3009 37323 3043
rect 37323 3009 37332 3043
rect 37280 3000 37332 3009
rect 37464 2975 37516 2984
rect 37464 2941 37473 2975
rect 37473 2941 37507 2975
rect 37507 2941 37516 2975
rect 37464 2932 37516 2941
rect 39672 3000 39724 3052
rect 40224 2932 40276 2984
rect 42156 2932 42208 2984
rect 44640 2932 44692 2984
rect 38016 2864 38068 2916
rect 41052 2864 41104 2916
rect 27896 2796 27948 2848
rect 31392 2796 31444 2848
rect 31760 2796 31812 2848
rect 34796 2796 34848 2848
rect 38660 2796 38712 2848
rect 43260 2864 43312 2916
rect 45468 2864 45520 2916
rect 46572 2864 46624 2916
rect 48228 2864 48280 2916
rect 49332 2864 49384 2916
rect 50988 2864 51040 2916
rect 52092 2864 52144 2916
rect 43812 2796 43864 2848
rect 46020 2796 46072 2848
rect 47400 2796 47452 2848
rect 48780 2796 48832 2848
rect 50160 2796 50212 2848
rect 51540 2796 51592 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 18144 2592 18196 2644
rect 22744 2592 22796 2644
rect 23848 2592 23900 2644
rect 25320 2592 25372 2644
rect 26608 2592 26660 2644
rect 28540 2592 28592 2644
rect 30380 2592 30432 2644
rect 30564 2592 30616 2644
rect 33140 2592 33192 2644
rect 33416 2592 33468 2644
rect 33876 2635 33928 2644
rect 33876 2601 33885 2635
rect 33885 2601 33919 2635
rect 33919 2601 33928 2635
rect 33876 2592 33928 2601
rect 34520 2635 34572 2644
rect 34520 2601 34529 2635
rect 34529 2601 34563 2635
rect 34563 2601 34572 2635
rect 34520 2592 34572 2601
rect 34704 2592 34756 2644
rect 36084 2592 36136 2644
rect 37464 2592 37516 2644
rect 37924 2592 37976 2644
rect 38660 2635 38712 2644
rect 38660 2601 38669 2635
rect 38669 2601 38703 2635
rect 38703 2601 38712 2635
rect 38660 2592 38712 2601
rect 39304 2635 39356 2644
rect 39304 2601 39313 2635
rect 39313 2601 39347 2635
rect 39347 2601 39356 2635
rect 39304 2592 39356 2601
rect 40040 2635 40092 2644
rect 40040 2601 40049 2635
rect 40049 2601 40083 2635
rect 40083 2601 40092 2635
rect 40040 2592 40092 2601
rect 47124 2592 47176 2644
rect 49884 2592 49936 2644
rect 10508 2524 10560 2576
rect 11888 2524 11940 2576
rect 13268 2524 13320 2576
rect 14648 2524 14700 2576
rect 17592 2524 17644 2576
rect 23112 2524 23164 2576
rect 25412 2524 25464 2576
rect 26792 2524 26844 2576
rect 29552 2524 29604 2576
rect 33600 2524 33652 2576
rect 35900 2524 35952 2576
rect 39396 2524 39448 2576
rect 42432 2524 42484 2576
rect 45192 2524 45244 2576
rect 47952 2524 48004 2576
rect 51264 2524 51316 2576
rect 16856 2456 16908 2508
rect 19340 2456 19392 2508
rect 7656 2388 7708 2440
rect 8208 2388 8260 2440
rect 8944 2388 8996 2440
rect 9680 2388 9732 2440
rect 11060 2388 11112 2440
rect 12440 2388 12492 2440
rect 13820 2388 13872 2440
rect 15476 2388 15528 2440
rect 19984 2388 20036 2440
rect 21364 2388 21416 2440
rect 24860 2456 24912 2508
rect 26516 2456 26568 2508
rect 30472 2456 30524 2508
rect 37188 2456 37240 2508
rect 41604 2456 41656 2508
rect 44088 2456 44140 2508
rect 46848 2456 46900 2508
rect 49608 2456 49660 2508
rect 52368 2456 52420 2508
rect 21456 2320 21508 2372
rect 23480 2431 23532 2440
rect 23480 2397 23489 2431
rect 23489 2397 23523 2431
rect 23523 2397 23532 2431
rect 23480 2388 23532 2397
rect 29644 2431 29696 2440
rect 29644 2397 29653 2431
rect 29653 2397 29687 2431
rect 29687 2397 29696 2431
rect 29644 2388 29696 2397
rect 32956 2388 33008 2440
rect 36728 2388 36780 2440
rect 24768 2320 24820 2372
rect 30656 2320 30708 2372
rect 37740 2320 37792 2372
rect 40776 2320 40828 2372
rect 42984 2388 43036 2440
rect 44364 2320 44416 2372
rect 45744 2320 45796 2372
rect 48504 2388 48556 2440
rect 50712 2320 50764 2372
rect 22744 2252 22796 2304
rect 25872 2252 25924 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 19984 2048 20036 2100
rect 23664 2048 23716 2100
rect 21364 1980 21416 2032
rect 25320 1980 25372 2032
rect 24860 1368 24912 1420
rect 25596 1368 25648 1420
<< metal2 >>
rect 3698 59200 3754 60000
rect 4158 59200 4214 60000
rect 4618 59200 4674 60000
rect 5078 59200 5134 60000
rect 5184 59214 5488 59242
rect 3712 57594 3740 59200
rect 3700 57588 3752 57594
rect 3700 57530 3752 57536
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4632 57050 4660 59200
rect 5092 59106 5120 59200
rect 5184 59106 5212 59214
rect 5092 59078 5212 59106
rect 5460 57610 5488 59214
rect 5538 59200 5594 60000
rect 5998 59200 6054 60000
rect 6458 59200 6514 60000
rect 6918 59200 6974 60000
rect 7378 59200 7434 60000
rect 7838 59200 7894 60000
rect 7944 59214 8248 59242
rect 5460 57594 5580 57610
rect 5460 57588 5592 57594
rect 5460 57582 5540 57588
rect 5540 57530 5592 57536
rect 6012 57050 6040 59200
rect 6366 57488 6422 57497
rect 6366 57423 6368 57432
rect 6420 57423 6422 57432
rect 6368 57394 6420 57400
rect 6472 57050 6500 59200
rect 7392 57458 7420 59200
rect 7852 59106 7880 59200
rect 7944 59106 7972 59214
rect 7852 59078 7972 59106
rect 8220 57882 8248 59214
rect 8298 59200 8354 60000
rect 8758 59200 8814 60000
rect 9218 59200 9274 60000
rect 9678 59200 9734 60000
rect 10138 59200 10194 60000
rect 10598 59200 10654 60000
rect 11058 59200 11114 60000
rect 11518 59200 11574 60000
rect 11978 59200 12034 60000
rect 12438 59200 12494 60000
rect 12898 59200 12954 60000
rect 13358 59200 13414 60000
rect 13818 59200 13874 60000
rect 14278 59200 14334 60000
rect 14738 59200 14794 60000
rect 15198 59200 15254 60000
rect 15658 59200 15714 60000
rect 16118 59200 16174 60000
rect 16578 59200 16634 60000
rect 17038 59200 17094 60000
rect 17498 59200 17554 60000
rect 17958 59200 18014 60000
rect 18418 59200 18474 60000
rect 18878 59200 18934 60000
rect 19338 59200 19394 60000
rect 19798 59200 19854 60000
rect 20258 59200 20314 60000
rect 20718 59200 20774 60000
rect 21178 59200 21234 60000
rect 21638 59200 21694 60000
rect 22098 59200 22154 60000
rect 22558 59200 22614 60000
rect 23018 59200 23074 60000
rect 23478 59200 23534 60000
rect 23938 59200 23994 60000
rect 24398 59200 24454 60000
rect 24858 59200 24914 60000
rect 25318 59200 25374 60000
rect 25778 59200 25834 60000
rect 26238 59200 26294 60000
rect 26698 59200 26754 60000
rect 27158 59200 27214 60000
rect 27264 59214 27568 59242
rect 8220 57854 8340 57882
rect 8312 57458 8340 57854
rect 7380 57452 7432 57458
rect 7380 57394 7432 57400
rect 8300 57452 8352 57458
rect 8300 57394 8352 57400
rect 8772 57050 8800 59200
rect 9232 57458 9260 59200
rect 9220 57452 9272 57458
rect 9220 57394 9272 57400
rect 10152 57050 10180 59200
rect 10612 57594 10640 59200
rect 10600 57588 10652 57594
rect 10600 57530 10652 57536
rect 11060 57316 11112 57322
rect 11060 57258 11112 57264
rect 4620 57044 4672 57050
rect 4620 56986 4672 56992
rect 6000 57044 6052 57050
rect 6000 56986 6052 56992
rect 6460 57044 6512 57050
rect 6460 56986 6512 56992
rect 8760 57044 8812 57050
rect 8760 56986 8812 56992
rect 10140 57044 10192 57050
rect 10140 56986 10192 56992
rect 11072 56914 11100 57258
rect 11532 57050 11560 59200
rect 11992 57594 12020 59200
rect 11980 57588 12032 57594
rect 11980 57530 12032 57536
rect 11888 57452 11940 57458
rect 11888 57394 11940 57400
rect 11900 57361 11928 57394
rect 11886 57352 11942 57361
rect 11886 57287 11942 57296
rect 12912 57050 12940 59200
rect 13268 57792 13320 57798
rect 13268 57734 13320 57740
rect 13280 57458 13308 57734
rect 13372 57594 13400 59200
rect 13360 57588 13412 57594
rect 13360 57530 13412 57536
rect 13268 57452 13320 57458
rect 13268 57394 13320 57400
rect 14292 57050 14320 59200
rect 14752 57594 14780 59200
rect 14740 57588 14792 57594
rect 14740 57530 14792 57536
rect 15672 57050 15700 59200
rect 16132 57594 16160 59200
rect 16120 57588 16172 57594
rect 16120 57530 16172 57536
rect 17052 57050 17080 59200
rect 17512 57594 17540 59200
rect 17500 57588 17552 57594
rect 17500 57530 17552 57536
rect 17408 57452 17460 57458
rect 17408 57394 17460 57400
rect 11520 57044 11572 57050
rect 11520 56986 11572 56992
rect 12900 57044 12952 57050
rect 12900 56986 12952 56992
rect 14280 57044 14332 57050
rect 14280 56986 14332 56992
rect 15660 57044 15712 57050
rect 15660 56986 15712 56992
rect 17040 57044 17092 57050
rect 17040 56986 17092 56992
rect 11060 56908 11112 56914
rect 11060 56850 11112 56856
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 17420 55894 17448 57394
rect 18432 57050 18460 59200
rect 18892 57594 18920 59200
rect 19812 58018 19840 59200
rect 19812 57990 20024 58018
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 18880 57588 18932 57594
rect 18880 57530 18932 57536
rect 19996 57050 20024 57990
rect 20168 57928 20220 57934
rect 20168 57870 20220 57876
rect 20180 57458 20208 57870
rect 20272 57594 20300 59200
rect 20260 57588 20312 57594
rect 20260 57530 20312 57536
rect 20168 57452 20220 57458
rect 20168 57394 20220 57400
rect 20720 57248 20772 57254
rect 20720 57190 20772 57196
rect 18420 57044 18472 57050
rect 18420 56986 18472 56992
rect 19984 57044 20036 57050
rect 19984 56986 20036 56992
rect 20732 56953 20760 57190
rect 21192 57050 21220 59200
rect 21652 57610 21680 59200
rect 21824 57860 21876 57866
rect 21824 57802 21876 57808
rect 21560 57594 21680 57610
rect 21548 57588 21680 57594
rect 21600 57582 21680 57588
rect 21548 57530 21600 57536
rect 21456 57520 21508 57526
rect 21732 57520 21784 57526
rect 21652 57480 21732 57508
rect 21652 57474 21680 57480
rect 21508 57468 21680 57474
rect 21456 57462 21680 57468
rect 21732 57462 21784 57468
rect 21468 57446 21680 57462
rect 21836 57458 21864 57802
rect 21824 57452 21876 57458
rect 21824 57394 21876 57400
rect 21916 57452 21968 57458
rect 21916 57394 21968 57400
rect 21928 57254 21956 57394
rect 22284 57384 22336 57390
rect 22284 57326 22336 57332
rect 21916 57248 21968 57254
rect 21916 57190 21968 57196
rect 22100 57248 22152 57254
rect 22100 57190 22152 57196
rect 21180 57044 21232 57050
rect 21180 56986 21232 56992
rect 20718 56944 20774 56953
rect 22112 56914 22140 57190
rect 22296 56982 22324 57326
rect 22284 56976 22336 56982
rect 22284 56918 22336 56924
rect 20718 56879 20774 56888
rect 22100 56908 22152 56914
rect 22100 56850 22152 56856
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 22572 56370 22600 59200
rect 23032 57050 23060 59200
rect 23756 57452 23808 57458
rect 23756 57394 23808 57400
rect 23664 57384 23716 57390
rect 23664 57326 23716 57332
rect 23020 57044 23072 57050
rect 23020 56986 23072 56992
rect 23204 56840 23256 56846
rect 23204 56782 23256 56788
rect 22560 56364 22612 56370
rect 22560 56306 22612 56312
rect 23216 56234 23244 56782
rect 23676 56302 23704 57326
rect 23768 56846 23796 57394
rect 23756 56840 23808 56846
rect 23756 56782 23808 56788
rect 23664 56296 23716 56302
rect 23664 56238 23716 56244
rect 23204 56228 23256 56234
rect 23204 56170 23256 56176
rect 23676 55962 23704 56238
rect 23768 55962 23796 56782
rect 23664 55956 23716 55962
rect 23664 55898 23716 55904
rect 23756 55956 23808 55962
rect 23756 55898 23808 55904
rect 17408 55888 17460 55894
rect 17408 55830 17460 55836
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 23952 55214 23980 59200
rect 24216 57792 24268 57798
rect 24216 57734 24268 57740
rect 24124 57452 24176 57458
rect 24124 57394 24176 57400
rect 24136 56846 24164 57394
rect 24228 57050 24256 57734
rect 24412 57594 24440 59200
rect 24492 57792 24544 57798
rect 24492 57734 24544 57740
rect 24400 57588 24452 57594
rect 24400 57530 24452 57536
rect 24308 57452 24360 57458
rect 24308 57394 24360 57400
rect 24216 57044 24268 57050
rect 24216 56986 24268 56992
rect 24124 56840 24176 56846
rect 24124 56782 24176 56788
rect 24032 56772 24084 56778
rect 24032 56714 24084 56720
rect 24044 56506 24072 56714
rect 24032 56500 24084 56506
rect 24032 56442 24084 56448
rect 24320 55758 24348 57394
rect 24504 56710 24532 57734
rect 25228 57452 25280 57458
rect 25228 57394 25280 57400
rect 25044 57316 25096 57322
rect 25044 57258 25096 57264
rect 25056 56710 25084 57258
rect 25240 56930 25268 57394
rect 25148 56902 25268 56930
rect 24492 56704 24544 56710
rect 24492 56646 24544 56652
rect 25044 56704 25096 56710
rect 25044 56646 25096 56652
rect 24504 56370 24532 56646
rect 24492 56364 24544 56370
rect 24492 56306 24544 56312
rect 25148 56302 25176 56902
rect 25136 56296 25188 56302
rect 25136 56238 25188 56244
rect 24308 55752 24360 55758
rect 24308 55694 24360 55700
rect 23940 55208 23992 55214
rect 23940 55150 23992 55156
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 25148 54874 25176 56238
rect 25332 55214 25360 59200
rect 25412 57928 25464 57934
rect 25412 57870 25464 57876
rect 25424 56914 25452 57870
rect 25504 57452 25556 57458
rect 25504 57394 25556 57400
rect 25412 56908 25464 56914
rect 25412 56850 25464 56856
rect 25424 55418 25452 56850
rect 25516 56846 25544 57394
rect 25596 57248 25648 57254
rect 25596 57190 25648 57196
rect 25504 56840 25556 56846
rect 25504 56782 25556 56788
rect 25504 56704 25556 56710
rect 25504 56646 25556 56652
rect 25516 56370 25544 56646
rect 25504 56364 25556 56370
rect 25504 56306 25556 56312
rect 25516 55865 25544 56306
rect 25502 55856 25558 55865
rect 25502 55791 25558 55800
rect 25412 55412 25464 55418
rect 25412 55354 25464 55360
rect 25320 55208 25372 55214
rect 25320 55150 25372 55156
rect 25136 54868 25188 54874
rect 25136 54810 25188 54816
rect 25608 54670 25636 57190
rect 25688 56160 25740 56166
rect 25688 56102 25740 56108
rect 25700 55282 25728 56102
rect 25792 55962 25820 59200
rect 26424 57860 26476 57866
rect 26424 57802 26476 57808
rect 26240 57384 26292 57390
rect 26240 57326 26292 57332
rect 25872 56908 25924 56914
rect 25872 56850 25924 56856
rect 25780 55956 25832 55962
rect 25780 55898 25832 55904
rect 25884 55758 25912 56850
rect 26252 56370 26280 57326
rect 26436 56914 26464 57802
rect 26424 56908 26476 56914
rect 26424 56850 26476 56856
rect 26516 56908 26568 56914
rect 26516 56850 26568 56856
rect 26240 56364 26292 56370
rect 26240 56306 26292 56312
rect 25872 55752 25924 55758
rect 25872 55694 25924 55700
rect 25688 55276 25740 55282
rect 25688 55218 25740 55224
rect 25884 54874 25912 55694
rect 26252 55282 26280 56306
rect 26240 55276 26292 55282
rect 26240 55218 26292 55224
rect 26252 54874 26280 55218
rect 26436 54874 26464 56850
rect 26528 55622 26556 56850
rect 26516 55616 26568 55622
rect 26516 55558 26568 55564
rect 25872 54868 25924 54874
rect 25872 54810 25924 54816
rect 26240 54868 26292 54874
rect 26240 54810 26292 54816
rect 26424 54868 26476 54874
rect 26424 54810 26476 54816
rect 25596 54664 25648 54670
rect 25596 54606 25648 54612
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 26252 54330 26280 54810
rect 26240 54324 26292 54330
rect 26240 54266 26292 54272
rect 26712 54194 26740 59200
rect 27172 59106 27200 59200
rect 27264 59106 27292 59214
rect 27172 59078 27292 59106
rect 27540 57769 27568 59214
rect 27618 59200 27674 60000
rect 27816 59214 28028 59242
rect 27712 57928 27764 57934
rect 27712 57870 27764 57876
rect 27526 57760 27582 57769
rect 27526 57695 27582 57704
rect 26976 57520 27028 57526
rect 26976 57462 27028 57468
rect 27160 57520 27212 57526
rect 27160 57462 27212 57468
rect 26884 57452 26936 57458
rect 26884 57394 26936 57400
rect 26896 56710 26924 57394
rect 26988 57050 27016 57462
rect 27068 57248 27120 57254
rect 27068 57190 27120 57196
rect 26976 57044 27028 57050
rect 26976 56986 27028 56992
rect 26884 56704 26936 56710
rect 26884 56646 26936 56652
rect 26896 56273 26924 56646
rect 26882 56264 26938 56273
rect 26882 56199 26938 56208
rect 27080 54670 27108 57190
rect 27172 56914 27200 57462
rect 27724 57458 27752 57870
rect 27712 57452 27764 57458
rect 27712 57394 27764 57400
rect 27620 57384 27672 57390
rect 27620 57326 27672 57332
rect 27710 57352 27766 57361
rect 27434 56944 27490 56953
rect 27160 56908 27212 56914
rect 27434 56879 27490 56888
rect 27160 56850 27212 56856
rect 27448 56846 27476 56879
rect 27344 56840 27396 56846
rect 27344 56782 27396 56788
rect 27436 56840 27488 56846
rect 27436 56782 27488 56788
rect 27526 56808 27582 56817
rect 27356 56370 27384 56782
rect 27526 56743 27528 56752
rect 27580 56743 27582 56752
rect 27528 56714 27580 56720
rect 27344 56364 27396 56370
rect 27344 56306 27396 56312
rect 27160 56160 27212 56166
rect 27160 56102 27212 56108
rect 27172 55826 27200 56102
rect 27160 55820 27212 55826
rect 27160 55762 27212 55768
rect 27356 55418 27384 56306
rect 27528 55820 27580 55826
rect 27528 55762 27580 55768
rect 27540 55690 27568 55762
rect 27528 55684 27580 55690
rect 27528 55626 27580 55632
rect 27344 55412 27396 55418
rect 27344 55354 27396 55360
rect 27632 55146 27660 57326
rect 27710 57287 27766 57296
rect 27724 57254 27752 57287
rect 27712 57248 27764 57254
rect 27712 57190 27764 57196
rect 27724 56914 27752 57190
rect 27712 56908 27764 56914
rect 27712 56850 27764 56856
rect 27710 56672 27766 56681
rect 27710 56607 27766 56616
rect 27724 56302 27752 56607
rect 27712 56296 27764 56302
rect 27712 56238 27764 56244
rect 27620 55140 27672 55146
rect 27620 55082 27672 55088
rect 27068 54664 27120 54670
rect 27068 54606 27120 54612
rect 26700 54188 26752 54194
rect 26700 54130 26752 54136
rect 27724 53990 27752 56238
rect 27816 55214 27844 59214
rect 28000 59106 28028 59214
rect 28078 59200 28134 60000
rect 28538 59200 28594 60000
rect 28644 59214 28948 59242
rect 28092 59106 28120 59200
rect 28000 59078 28120 59106
rect 28552 59106 28580 59200
rect 28644 59106 28672 59214
rect 28552 59078 28672 59106
rect 28080 57860 28132 57866
rect 28080 57802 28132 57808
rect 27986 57488 28042 57497
rect 27896 57452 27948 57458
rect 27986 57423 28042 57432
rect 27896 57394 27948 57400
rect 27908 56438 27936 57394
rect 28000 56982 28028 57423
rect 28092 57050 28120 57802
rect 28170 57760 28226 57769
rect 28170 57695 28226 57704
rect 28184 57526 28212 57695
rect 28920 57610 28948 59214
rect 28998 59200 29054 60000
rect 29458 59200 29514 60000
rect 29564 59214 29776 59242
rect 29012 57746 29040 59200
rect 29472 59106 29500 59200
rect 29564 59106 29592 59214
rect 29472 59078 29592 59106
rect 29012 57718 29132 57746
rect 28920 57594 29040 57610
rect 28920 57588 29052 57594
rect 28920 57582 29000 57588
rect 29000 57530 29052 57536
rect 28172 57520 28224 57526
rect 28172 57462 28224 57468
rect 28172 57384 28224 57390
rect 28172 57326 28224 57332
rect 28184 57050 28212 57326
rect 28264 57316 28316 57322
rect 28264 57258 28316 57264
rect 28908 57316 28960 57322
rect 28908 57258 28960 57264
rect 28080 57044 28132 57050
rect 28080 56986 28132 56992
rect 28172 57044 28224 57050
rect 28172 56986 28224 56992
rect 27988 56976 28040 56982
rect 27988 56918 28040 56924
rect 28172 56840 28224 56846
rect 28172 56782 28224 56788
rect 28080 56772 28132 56778
rect 28080 56714 28132 56720
rect 27896 56432 27948 56438
rect 27896 56374 27948 56380
rect 27988 56296 28040 56302
rect 27988 56238 28040 56244
rect 28000 55690 28028 56238
rect 27988 55684 28040 55690
rect 27988 55626 28040 55632
rect 27804 55208 27856 55214
rect 27804 55150 27856 55156
rect 27712 53984 27764 53990
rect 27712 53926 27764 53932
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 27724 8090 27752 53926
rect 28092 53786 28120 56714
rect 28184 56506 28212 56782
rect 28172 56500 28224 56506
rect 28172 56442 28224 56448
rect 28276 56370 28304 57258
rect 28920 56982 28948 57258
rect 28448 56976 28500 56982
rect 28448 56918 28500 56924
rect 28908 56976 28960 56982
rect 28908 56918 28960 56924
rect 28264 56364 28316 56370
rect 28264 56306 28316 56312
rect 28276 55894 28304 56306
rect 28264 55888 28316 55894
rect 28264 55830 28316 55836
rect 28264 55616 28316 55622
rect 28264 55558 28316 55564
rect 28276 55146 28304 55558
rect 28264 55140 28316 55146
rect 28264 55082 28316 55088
rect 28460 54738 28488 56918
rect 28540 56772 28592 56778
rect 28540 56714 28592 56720
rect 28448 54732 28500 54738
rect 28448 54674 28500 54680
rect 28552 54670 28580 56714
rect 28632 56432 28684 56438
rect 28632 56374 28684 56380
rect 28644 55894 28672 56374
rect 29000 56160 29052 56166
rect 29000 56102 29052 56108
rect 29012 55962 29040 56102
rect 29000 55956 29052 55962
rect 29000 55898 29052 55904
rect 28632 55888 28684 55894
rect 28632 55830 28684 55836
rect 28816 55752 28868 55758
rect 28816 55694 28868 55700
rect 28908 55752 28960 55758
rect 28908 55694 28960 55700
rect 28828 55214 28856 55694
rect 28920 55622 28948 55694
rect 28908 55616 28960 55622
rect 28908 55558 28960 55564
rect 29104 55298 29132 57718
rect 29644 57588 29696 57594
rect 29644 57530 29696 57536
rect 29460 57452 29512 57458
rect 29460 57394 29512 57400
rect 29196 57310 29408 57338
rect 29196 56914 29224 57310
rect 29380 57254 29408 57310
rect 29276 57248 29328 57254
rect 29276 57190 29328 57196
rect 29368 57248 29420 57254
rect 29368 57190 29420 57196
rect 29184 56908 29236 56914
rect 29184 56850 29236 56856
rect 29288 56846 29316 57190
rect 29368 56976 29420 56982
rect 29368 56918 29420 56924
rect 29380 56846 29408 56918
rect 29276 56840 29328 56846
rect 29276 56782 29328 56788
rect 29368 56840 29420 56846
rect 29368 56782 29420 56788
rect 29288 56352 29316 56782
rect 29472 56710 29500 57394
rect 29552 56976 29604 56982
rect 29552 56918 29604 56924
rect 29460 56704 29512 56710
rect 29460 56646 29512 56652
rect 29196 56324 29316 56352
rect 29366 56400 29422 56409
rect 29472 56370 29500 56646
rect 29366 56335 29368 56344
rect 29196 55826 29224 56324
rect 29420 56335 29422 56344
rect 29460 56364 29512 56370
rect 29368 56306 29420 56312
rect 29460 56306 29512 56312
rect 29564 56250 29592 56918
rect 29276 56228 29328 56234
rect 29276 56170 29328 56176
rect 29472 56222 29592 56250
rect 29184 55820 29236 55826
rect 29184 55762 29236 55768
rect 28920 55270 29132 55298
rect 29184 55276 29236 55282
rect 28816 55208 28868 55214
rect 28816 55150 28868 55156
rect 28724 55072 28776 55078
rect 28724 55014 28776 55020
rect 28736 54738 28764 55014
rect 28724 54732 28776 54738
rect 28724 54674 28776 54680
rect 28540 54664 28592 54670
rect 28540 54606 28592 54612
rect 28920 54194 28948 55270
rect 29184 55218 29236 55224
rect 29000 54664 29052 54670
rect 29000 54606 29052 54612
rect 28908 54188 28960 54194
rect 28908 54130 28960 54136
rect 28920 53786 28948 54130
rect 29012 53786 29040 54606
rect 28080 53780 28132 53786
rect 28080 53722 28132 53728
rect 28908 53780 28960 53786
rect 28908 53722 28960 53728
rect 29000 53780 29052 53786
rect 29000 53722 29052 53728
rect 29196 53582 29224 55218
rect 29288 54874 29316 56170
rect 29368 55276 29420 55282
rect 29368 55218 29420 55224
rect 29276 54868 29328 54874
rect 29276 54810 29328 54816
rect 29380 54330 29408 55218
rect 29472 54806 29500 56222
rect 29656 55758 29684 57530
rect 29644 55752 29696 55758
rect 29644 55694 29696 55700
rect 29460 54800 29512 54806
rect 29460 54742 29512 54748
rect 29368 54324 29420 54330
rect 29368 54266 29420 54272
rect 29184 53576 29236 53582
rect 29184 53518 29236 53524
rect 29380 53446 29408 54266
rect 29472 54262 29500 54742
rect 29460 54256 29512 54262
rect 29460 54198 29512 54204
rect 29748 53786 29776 59214
rect 29918 59200 29974 60000
rect 30378 59200 30434 60000
rect 30838 59200 30894 60000
rect 31298 59200 31354 60000
rect 31758 59200 31814 60000
rect 32218 59200 32274 60000
rect 32678 59200 32734 60000
rect 33138 59200 33194 60000
rect 33244 59214 33548 59242
rect 29828 56840 29880 56846
rect 29828 56782 29880 56788
rect 29840 56681 29868 56782
rect 29826 56672 29882 56681
rect 29826 56607 29882 56616
rect 29826 56536 29882 56545
rect 29826 56471 29882 56480
rect 29840 56370 29868 56471
rect 29828 56364 29880 56370
rect 29828 56306 29880 56312
rect 29828 55616 29880 55622
rect 29828 55558 29880 55564
rect 29840 55457 29868 55558
rect 29826 55448 29882 55457
rect 29826 55383 29882 55392
rect 29932 54874 29960 59200
rect 30392 57610 30420 59200
rect 30300 57594 30420 57610
rect 30288 57588 30420 57594
rect 30340 57582 30420 57588
rect 30656 57588 30708 57594
rect 30288 57530 30340 57536
rect 30656 57530 30708 57536
rect 30668 57254 30696 57530
rect 30656 57248 30708 57254
rect 30656 57190 30708 57196
rect 30010 56808 30066 56817
rect 30010 56743 30066 56752
rect 30024 56710 30052 56743
rect 30012 56704 30064 56710
rect 30012 56646 30064 56652
rect 30472 56500 30524 56506
rect 30472 56442 30524 56448
rect 30196 56364 30248 56370
rect 30196 56306 30248 56312
rect 30104 56160 30156 56166
rect 30104 56102 30156 56108
rect 30012 55616 30064 55622
rect 30012 55558 30064 55564
rect 30024 55418 30052 55558
rect 30116 55418 30144 56102
rect 30208 55962 30236 56306
rect 30484 56302 30512 56442
rect 30748 56432 30800 56438
rect 30748 56374 30800 56380
rect 30472 56296 30524 56302
rect 30472 56238 30524 56244
rect 30196 55956 30248 55962
rect 30196 55898 30248 55904
rect 30208 55690 30236 55898
rect 30380 55820 30432 55826
rect 30380 55762 30432 55768
rect 30288 55752 30340 55758
rect 30288 55694 30340 55700
rect 30196 55684 30248 55690
rect 30196 55626 30248 55632
rect 30300 55418 30328 55694
rect 30012 55412 30064 55418
rect 30012 55354 30064 55360
rect 30104 55412 30156 55418
rect 30104 55354 30156 55360
rect 30288 55412 30340 55418
rect 30288 55354 30340 55360
rect 30392 55282 30420 55762
rect 30472 55344 30524 55350
rect 30472 55286 30524 55292
rect 30012 55276 30064 55282
rect 30012 55218 30064 55224
rect 30380 55276 30432 55282
rect 30380 55218 30432 55224
rect 29920 54868 29972 54874
rect 29920 54810 29972 54816
rect 30024 54330 30052 55218
rect 30288 55208 30340 55214
rect 30288 55150 30340 55156
rect 30196 54732 30248 54738
rect 30196 54674 30248 54680
rect 30012 54324 30064 54330
rect 30012 54266 30064 54272
rect 29736 53780 29788 53786
rect 29736 53722 29788 53728
rect 30024 53582 30052 54266
rect 30208 54194 30236 54674
rect 30300 54330 30328 55150
rect 30484 54874 30512 55286
rect 30472 54868 30524 54874
rect 30472 54810 30524 54816
rect 30380 54596 30432 54602
rect 30380 54538 30432 54544
rect 30288 54324 30340 54330
rect 30288 54266 30340 54272
rect 30392 54194 30420 54538
rect 30760 54262 30788 56374
rect 30852 56370 30880 59200
rect 31024 57248 31076 57254
rect 31024 57190 31076 57196
rect 31036 56846 31064 57190
rect 31024 56840 31076 56846
rect 31024 56782 31076 56788
rect 30840 56364 30892 56370
rect 30840 56306 30892 56312
rect 31036 55826 31064 56782
rect 31024 55820 31076 55826
rect 31024 55762 31076 55768
rect 30932 55684 30984 55690
rect 30932 55626 30984 55632
rect 30944 55418 30972 55626
rect 30932 55412 30984 55418
rect 30932 55354 30984 55360
rect 30748 54256 30800 54262
rect 30748 54198 30800 54204
rect 31036 54194 31064 55762
rect 31312 54874 31340 59200
rect 31772 57458 31800 59200
rect 31760 57452 31812 57458
rect 31760 57394 31812 57400
rect 31772 56930 31800 57394
rect 32232 57254 32260 59200
rect 32404 57384 32456 57390
rect 32404 57326 32456 57332
rect 32220 57248 32272 57254
rect 32220 57190 32272 57196
rect 31772 56902 31984 56930
rect 31760 56840 31812 56846
rect 31812 56788 31892 56794
rect 31760 56782 31892 56788
rect 31772 56766 31892 56782
rect 31760 56704 31812 56710
rect 31760 56646 31812 56652
rect 31772 56370 31800 56646
rect 31864 56506 31892 56766
rect 31852 56500 31904 56506
rect 31852 56442 31904 56448
rect 31760 56364 31812 56370
rect 31760 56306 31812 56312
rect 31852 56160 31904 56166
rect 31852 56102 31904 56108
rect 31864 55078 31892 56102
rect 31852 55072 31904 55078
rect 31852 55014 31904 55020
rect 31300 54868 31352 54874
rect 31300 54810 31352 54816
rect 30196 54188 30248 54194
rect 30196 54130 30248 54136
rect 30380 54188 30432 54194
rect 30380 54130 30432 54136
rect 31024 54188 31076 54194
rect 31024 54130 31076 54136
rect 31036 53786 31064 54130
rect 31864 54058 31892 55014
rect 31852 54052 31904 54058
rect 31852 53994 31904 54000
rect 31956 53786 31984 56902
rect 32220 56772 32272 56778
rect 32220 56714 32272 56720
rect 32036 56704 32088 56710
rect 32036 56646 32088 56652
rect 32048 56166 32076 56646
rect 32232 56370 32260 56714
rect 32220 56364 32272 56370
rect 32220 56306 32272 56312
rect 32036 56160 32088 56166
rect 32036 56102 32088 56108
rect 32128 55752 32180 55758
rect 32128 55694 32180 55700
rect 32140 55350 32168 55694
rect 32128 55344 32180 55350
rect 32128 55286 32180 55292
rect 32232 55282 32260 56306
rect 32416 55758 32444 57326
rect 32692 57202 32720 59200
rect 33152 59106 33180 59200
rect 33244 59106 33272 59214
rect 33152 59078 33272 59106
rect 32956 57520 33008 57526
rect 32956 57462 33008 57468
rect 32692 57174 32812 57202
rect 32680 57044 32732 57050
rect 32680 56986 32732 56992
rect 32692 56506 32720 56986
rect 32680 56500 32732 56506
rect 32680 56442 32732 56448
rect 32404 55752 32456 55758
rect 32404 55694 32456 55700
rect 32220 55276 32272 55282
rect 32220 55218 32272 55224
rect 32312 55072 32364 55078
rect 32312 55014 32364 55020
rect 32324 54738 32352 55014
rect 32312 54732 32364 54738
rect 32312 54674 32364 54680
rect 32324 54176 32352 54674
rect 32416 54602 32444 55694
rect 32784 55282 32812 57174
rect 32968 55457 32996 57462
rect 33416 57316 33468 57322
rect 33416 57258 33468 57264
rect 33428 56846 33456 57258
rect 33416 56840 33468 56846
rect 33416 56782 33468 56788
rect 33232 56704 33284 56710
rect 33232 56646 33284 56652
rect 33244 56370 33272 56646
rect 33232 56364 33284 56370
rect 33232 56306 33284 56312
rect 33140 56296 33192 56302
rect 33140 56238 33192 56244
rect 33048 56160 33100 56166
rect 33048 56102 33100 56108
rect 32954 55448 33010 55457
rect 32954 55383 33010 55392
rect 32772 55276 32824 55282
rect 32772 55218 32824 55224
rect 32772 55072 32824 55078
rect 32772 55014 32824 55020
rect 32784 54670 32812 55014
rect 32772 54664 32824 54670
rect 32772 54606 32824 54612
rect 32404 54596 32456 54602
rect 32404 54538 32456 54544
rect 32968 54194 32996 55383
rect 33060 54806 33088 56102
rect 33152 55622 33180 56238
rect 33428 55758 33456 56782
rect 33416 55752 33468 55758
rect 33416 55694 33468 55700
rect 33140 55616 33192 55622
rect 33140 55558 33192 55564
rect 33140 55276 33192 55282
rect 33140 55218 33192 55224
rect 33048 54800 33100 54806
rect 33048 54742 33100 54748
rect 33152 54330 33180 55218
rect 33416 55072 33468 55078
rect 33416 55014 33468 55020
rect 33324 54528 33376 54534
rect 33324 54470 33376 54476
rect 33140 54324 33192 54330
rect 33140 54266 33192 54272
rect 33232 54256 33284 54262
rect 33232 54198 33284 54204
rect 32404 54188 32456 54194
rect 32324 54148 32404 54176
rect 32404 54130 32456 54136
rect 32956 54188 33008 54194
rect 32956 54130 33008 54136
rect 33140 54188 33192 54194
rect 33140 54130 33192 54136
rect 31024 53780 31076 53786
rect 31024 53722 31076 53728
rect 31944 53780 31996 53786
rect 31944 53722 31996 53728
rect 30012 53576 30064 53582
rect 30012 53518 30064 53524
rect 29368 53440 29420 53446
rect 29368 53382 29420 53388
rect 31036 53242 31064 53722
rect 32588 53644 32640 53650
rect 32588 53586 32640 53592
rect 32600 53242 32628 53586
rect 33152 53582 33180 54130
rect 33244 53786 33272 54198
rect 33336 54194 33364 54470
rect 33324 54188 33376 54194
rect 33324 54130 33376 54136
rect 33232 53780 33284 53786
rect 33232 53722 33284 53728
rect 33140 53576 33192 53582
rect 33140 53518 33192 53524
rect 33336 53514 33364 54130
rect 33428 54126 33456 55014
rect 33520 54194 33548 59214
rect 33598 59200 33654 60000
rect 34058 59200 34114 60000
rect 34518 59200 34574 60000
rect 34978 59200 35034 60000
rect 35084 59214 35388 59242
rect 33612 55282 33640 59200
rect 33692 57452 33744 57458
rect 33692 57394 33744 57400
rect 33784 57452 33836 57458
rect 33784 57394 33836 57400
rect 33704 56234 33732 57394
rect 33796 56846 33824 57394
rect 33784 56840 33836 56846
rect 33784 56782 33836 56788
rect 33692 56228 33744 56234
rect 33692 56170 33744 56176
rect 33600 55276 33652 55282
rect 33600 55218 33652 55224
rect 33704 54330 33732 56170
rect 33876 56160 33928 56166
rect 33876 56102 33928 56108
rect 33968 56160 34020 56166
rect 33968 56102 34020 56108
rect 33888 55078 33916 56102
rect 33980 55894 34008 56102
rect 34072 55894 34100 59200
rect 34336 57248 34388 57254
rect 34336 57190 34388 57196
rect 34348 56914 34376 57190
rect 34336 56908 34388 56914
rect 34336 56850 34388 56856
rect 34428 56840 34480 56846
rect 34428 56782 34480 56788
rect 34440 55962 34468 56782
rect 34532 56506 34560 59200
rect 34992 59106 35020 59200
rect 35084 59106 35112 59214
rect 34992 59078 35112 59106
rect 34704 57928 34756 57934
rect 34704 57870 34756 57876
rect 34612 57316 34664 57322
rect 34612 57258 34664 57264
rect 34624 56846 34652 57258
rect 34612 56840 34664 56846
rect 34612 56782 34664 56788
rect 34716 56794 34744 57870
rect 34796 57452 34848 57458
rect 34796 57394 34848 57400
rect 34808 56982 34836 57394
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 34796 56976 34848 56982
rect 34796 56918 34848 56924
rect 34900 56846 34928 56877
rect 34888 56840 34940 56846
rect 34716 56788 34888 56794
rect 34716 56782 34940 56788
rect 34624 56692 34652 56782
rect 34716 56766 34928 56782
rect 34624 56664 34744 56692
rect 34520 56500 34572 56506
rect 34520 56442 34572 56448
rect 34716 56438 34744 56664
rect 34796 56500 34848 56506
rect 34796 56442 34848 56448
rect 34704 56432 34756 56438
rect 34704 56374 34756 56380
rect 34612 56364 34664 56370
rect 34612 56306 34664 56312
rect 34428 55956 34480 55962
rect 34428 55898 34480 55904
rect 33968 55888 34020 55894
rect 33968 55830 34020 55836
rect 34060 55888 34112 55894
rect 34060 55830 34112 55836
rect 34624 55826 34652 56306
rect 34612 55820 34664 55826
rect 34612 55762 34664 55768
rect 34624 55418 34652 55762
rect 34716 55758 34744 56374
rect 34704 55752 34756 55758
rect 34704 55694 34756 55700
rect 34612 55412 34664 55418
rect 34612 55354 34664 55360
rect 33876 55072 33928 55078
rect 33876 55014 33928 55020
rect 33888 54738 33916 55014
rect 33876 54732 33928 54738
rect 33876 54674 33928 54680
rect 33692 54324 33744 54330
rect 33692 54266 33744 54272
rect 33508 54188 33560 54194
rect 33508 54130 33560 54136
rect 33968 54188 34020 54194
rect 33968 54130 34020 54136
rect 33416 54120 33468 54126
rect 33416 54062 33468 54068
rect 33428 53718 33456 54062
rect 33980 53786 34008 54130
rect 34808 53786 34836 56442
rect 34900 56438 34928 56766
rect 34888 56432 34940 56438
rect 34888 56374 34940 56380
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34888 54800 34940 54806
rect 34888 54742 34940 54748
rect 34900 54194 34928 54742
rect 35360 54194 35388 59214
rect 35438 59200 35494 60000
rect 35898 59200 35954 60000
rect 36358 59200 36414 60000
rect 36818 59200 36874 60000
rect 37278 59200 37334 60000
rect 37738 59200 37794 60000
rect 38198 59200 38254 60000
rect 38658 59200 38714 60000
rect 39118 59200 39174 60000
rect 39578 59200 39634 60000
rect 40038 59200 40094 60000
rect 40498 59200 40554 60000
rect 40958 59200 41014 60000
rect 41418 59200 41474 60000
rect 41524 59214 41736 59242
rect 35452 55350 35480 59200
rect 35532 57588 35584 57594
rect 35532 57530 35584 57536
rect 35544 56506 35572 57530
rect 35624 57520 35676 57526
rect 35624 57462 35676 57468
rect 35532 56500 35584 56506
rect 35532 56442 35584 56448
rect 35532 56364 35584 56370
rect 35532 56306 35584 56312
rect 35440 55344 35492 55350
rect 35440 55286 35492 55292
rect 34888 54188 34940 54194
rect 34888 54130 34940 54136
rect 35348 54188 35400 54194
rect 35348 54130 35400 54136
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 33968 53780 34020 53786
rect 33968 53722 34020 53728
rect 34796 53780 34848 53786
rect 34796 53722 34848 53728
rect 33416 53712 33468 53718
rect 33416 53654 33468 53660
rect 33324 53508 33376 53514
rect 33324 53450 33376 53456
rect 31024 53236 31076 53242
rect 31024 53178 31076 53184
rect 32588 53236 32640 53242
rect 32588 53178 32640 53184
rect 35544 53174 35572 56306
rect 35636 55418 35664 57462
rect 35912 57390 35940 59200
rect 36176 57860 36228 57866
rect 36176 57802 36228 57808
rect 35900 57384 35952 57390
rect 35900 57326 35952 57332
rect 35624 55412 35676 55418
rect 35624 55354 35676 55360
rect 35636 54670 35664 55354
rect 35716 55072 35768 55078
rect 35716 55014 35768 55020
rect 35728 54670 35756 55014
rect 35624 54664 35676 54670
rect 35624 54606 35676 54612
rect 35716 54664 35768 54670
rect 35716 54606 35768 54612
rect 35728 54126 35756 54606
rect 35716 54120 35768 54126
rect 35716 54062 35768 54068
rect 35912 53718 35940 57326
rect 36084 56704 36136 56710
rect 36084 56646 36136 56652
rect 36096 56545 36124 56646
rect 36082 56536 36138 56545
rect 36188 56506 36216 57802
rect 36268 57452 36320 57458
rect 36268 57394 36320 57400
rect 36082 56471 36138 56480
rect 36176 56500 36228 56506
rect 36176 56442 36228 56448
rect 36176 56160 36228 56166
rect 36176 56102 36228 56108
rect 35992 55888 36044 55894
rect 35992 55830 36044 55836
rect 36004 55146 36032 55830
rect 36084 55820 36136 55826
rect 36084 55762 36136 55768
rect 35992 55140 36044 55146
rect 35992 55082 36044 55088
rect 36096 53786 36124 55762
rect 36188 55622 36216 56102
rect 36176 55616 36228 55622
rect 36176 55558 36228 55564
rect 36188 55282 36216 55558
rect 36176 55276 36228 55282
rect 36176 55218 36228 55224
rect 36188 54670 36216 55218
rect 36280 55214 36308 57394
rect 36268 55208 36320 55214
rect 36268 55150 36320 55156
rect 36280 54874 36308 55150
rect 36372 54874 36400 59200
rect 36452 57248 36504 57254
rect 36452 57190 36504 57196
rect 36464 56778 36492 57190
rect 36452 56772 36504 56778
rect 36452 56714 36504 56720
rect 36464 55690 36492 56714
rect 36452 55684 36504 55690
rect 36452 55626 36504 55632
rect 36268 54868 36320 54874
rect 36268 54810 36320 54816
rect 36360 54868 36412 54874
rect 36360 54810 36412 54816
rect 36176 54664 36228 54670
rect 36176 54606 36228 54612
rect 36188 54262 36216 54606
rect 36464 54330 36492 55626
rect 36832 55282 36860 59200
rect 37292 57390 37320 59200
rect 37280 57384 37332 57390
rect 37280 57326 37332 57332
rect 37464 57384 37516 57390
rect 37464 57326 37516 57332
rect 37372 57044 37424 57050
rect 37372 56986 37424 56992
rect 37280 56840 37332 56846
rect 37280 56782 37332 56788
rect 37292 56506 37320 56782
rect 37280 56500 37332 56506
rect 37280 56442 37332 56448
rect 37384 56409 37412 56986
rect 37370 56400 37426 56409
rect 37370 56335 37426 56344
rect 37002 55992 37058 56001
rect 37002 55927 37058 55936
rect 37016 55758 37044 55927
rect 37004 55752 37056 55758
rect 37004 55694 37056 55700
rect 36820 55276 36872 55282
rect 36820 55218 36872 55224
rect 37280 55276 37332 55282
rect 37280 55218 37332 55224
rect 36452 54324 36504 54330
rect 36452 54266 36504 54272
rect 36176 54256 36228 54262
rect 36176 54198 36228 54204
rect 36084 53780 36136 53786
rect 36084 53722 36136 53728
rect 35900 53712 35952 53718
rect 35900 53654 35952 53660
rect 35992 53644 36044 53650
rect 35992 53586 36044 53592
rect 35532 53168 35584 53174
rect 35532 53110 35584 53116
rect 34796 53032 34848 53038
rect 34796 52974 34848 52980
rect 34808 45554 34836 52974
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 36004 52698 36032 53586
rect 36096 53242 36124 53722
rect 36464 53650 36492 54266
rect 37292 54194 37320 55218
rect 37280 54188 37332 54194
rect 37280 54130 37332 54136
rect 37476 53786 37504 57326
rect 37648 56364 37700 56370
rect 37648 56306 37700 56312
rect 37660 55758 37688 56306
rect 37648 55752 37700 55758
rect 37648 55694 37700 55700
rect 37752 54194 37780 59200
rect 37832 56908 37884 56914
rect 37832 56850 37884 56856
rect 37844 56438 37872 56850
rect 37832 56432 37884 56438
rect 37832 56374 37884 56380
rect 38108 56228 38160 56234
rect 38108 56170 38160 56176
rect 37830 55992 37886 56001
rect 37830 55927 37886 55936
rect 37844 54670 37872 55927
rect 38016 55888 38068 55894
rect 38016 55830 38068 55836
rect 37924 55684 37976 55690
rect 37924 55626 37976 55632
rect 37936 55418 37964 55626
rect 38028 55457 38056 55830
rect 38014 55448 38070 55457
rect 37924 55412 37976 55418
rect 38014 55383 38070 55392
rect 37924 55354 37976 55360
rect 38028 54670 38056 55383
rect 38120 54874 38148 56170
rect 38108 54868 38160 54874
rect 38108 54810 38160 54816
rect 37832 54664 37884 54670
rect 37832 54606 37884 54612
rect 38016 54664 38068 54670
rect 38016 54606 38068 54612
rect 38212 54194 38240 59200
rect 38672 57458 38700 59200
rect 39132 57934 39160 59200
rect 39120 57928 39172 57934
rect 39120 57870 39172 57876
rect 38660 57452 38712 57458
rect 38660 57394 38712 57400
rect 38844 56840 38896 56846
rect 38844 56782 38896 56788
rect 38936 56840 38988 56846
rect 38936 56782 38988 56788
rect 38856 56370 38884 56782
rect 38844 56364 38896 56370
rect 38844 56306 38896 56312
rect 38568 56296 38620 56302
rect 38568 56238 38620 56244
rect 38292 55888 38344 55894
rect 38292 55830 38344 55836
rect 38304 55758 38332 55830
rect 38580 55826 38608 56238
rect 38948 56234 38976 56782
rect 39212 56364 39264 56370
rect 39212 56306 39264 56312
rect 38936 56228 38988 56234
rect 38936 56170 38988 56176
rect 39224 55962 39252 56306
rect 39212 55956 39264 55962
rect 39212 55898 39264 55904
rect 38568 55820 38620 55826
rect 38568 55762 38620 55768
rect 38292 55752 38344 55758
rect 38292 55694 38344 55700
rect 38936 55752 38988 55758
rect 38936 55694 38988 55700
rect 39488 55752 39540 55758
rect 39488 55694 39540 55700
rect 38948 55622 38976 55694
rect 38936 55616 38988 55622
rect 38936 55558 38988 55564
rect 38752 55344 38804 55350
rect 38752 55286 38804 55292
rect 38764 55214 38792 55286
rect 38752 55208 38804 55214
rect 38752 55150 38804 55156
rect 38764 54670 38792 55150
rect 38948 54874 38976 55558
rect 39028 55140 39080 55146
rect 39028 55082 39080 55088
rect 38936 54868 38988 54874
rect 38936 54810 38988 54816
rect 39040 54670 39068 55082
rect 39500 54670 39528 55694
rect 38752 54664 38804 54670
rect 38752 54606 38804 54612
rect 39028 54664 39080 54670
rect 39028 54606 39080 54612
rect 39488 54664 39540 54670
rect 39488 54606 39540 54612
rect 39592 54194 39620 59200
rect 39948 57792 40000 57798
rect 39948 57734 40000 57740
rect 39960 57594 39988 57734
rect 39948 57588 40000 57594
rect 39948 57530 40000 57536
rect 39856 57452 39908 57458
rect 39856 57394 39908 57400
rect 39764 56976 39816 56982
rect 39764 56918 39816 56924
rect 39776 56370 39804 56918
rect 39764 56364 39816 56370
rect 39764 56306 39816 56312
rect 39672 55072 39724 55078
rect 39672 55014 39724 55020
rect 39684 54670 39712 55014
rect 39776 54806 39804 56306
rect 39764 54800 39816 54806
rect 39764 54742 39816 54748
rect 39672 54664 39724 54670
rect 39672 54606 39724 54612
rect 39684 54330 39712 54606
rect 39672 54324 39724 54330
rect 39672 54266 39724 54272
rect 37740 54188 37792 54194
rect 37740 54130 37792 54136
rect 38200 54188 38252 54194
rect 38200 54130 38252 54136
rect 39580 54188 39632 54194
rect 39580 54130 39632 54136
rect 37464 53780 37516 53786
rect 37464 53722 37516 53728
rect 39868 53718 39896 57394
rect 40052 56953 40080 59200
rect 40132 57860 40184 57866
rect 40132 57802 40184 57808
rect 40144 57254 40172 57802
rect 40512 57798 40540 59200
rect 40500 57792 40552 57798
rect 40500 57734 40552 57740
rect 40224 57520 40276 57526
rect 40224 57462 40276 57468
rect 40132 57248 40184 57254
rect 40132 57190 40184 57196
rect 40038 56944 40094 56953
rect 40038 56879 40094 56888
rect 40144 56846 40172 57190
rect 40236 56846 40264 57462
rect 40316 57384 40368 57390
rect 40500 57384 40552 57390
rect 40368 57344 40448 57372
rect 40316 57326 40368 57332
rect 40420 56982 40448 57344
rect 40500 57326 40552 57332
rect 40408 56976 40460 56982
rect 40408 56918 40460 56924
rect 40132 56840 40184 56846
rect 40132 56782 40184 56788
rect 40224 56840 40276 56846
rect 40224 56782 40276 56788
rect 40132 56364 40184 56370
rect 40132 56306 40184 56312
rect 40040 56296 40092 56302
rect 40040 56238 40092 56244
rect 40052 54058 40080 56238
rect 40144 54874 40172 56306
rect 40236 55826 40264 56782
rect 40316 56704 40368 56710
rect 40316 56646 40368 56652
rect 40224 55820 40276 55826
rect 40224 55762 40276 55768
rect 40236 55282 40264 55762
rect 40328 55758 40356 56646
rect 40420 56302 40448 56918
rect 40408 56296 40460 56302
rect 40408 56238 40460 56244
rect 40316 55752 40368 55758
rect 40316 55694 40368 55700
rect 40224 55276 40276 55282
rect 40224 55218 40276 55224
rect 40132 54868 40184 54874
rect 40132 54810 40184 54816
rect 40316 54732 40368 54738
rect 40316 54674 40368 54680
rect 40328 54194 40356 54674
rect 40420 54262 40448 56238
rect 40512 55962 40540 57326
rect 40592 57316 40644 57322
rect 40592 57258 40644 57264
rect 40604 56710 40632 57258
rect 40776 57248 40828 57254
rect 40776 57190 40828 57196
rect 40592 56704 40644 56710
rect 40590 56672 40592 56681
rect 40644 56672 40646 56681
rect 40590 56607 40646 56616
rect 40500 55956 40552 55962
rect 40500 55898 40552 55904
rect 40604 55894 40632 56607
rect 40788 56438 40816 57190
rect 40972 56522 41000 59200
rect 41432 59106 41460 59200
rect 41524 59106 41552 59214
rect 41432 59078 41552 59106
rect 41328 56704 41380 56710
rect 41328 56646 41380 56652
rect 40972 56494 41092 56522
rect 40776 56432 40828 56438
rect 40776 56374 40828 56380
rect 40960 56364 41012 56370
rect 40960 56306 41012 56312
rect 40682 56264 40738 56273
rect 40682 56199 40684 56208
rect 40736 56199 40738 56208
rect 40684 56170 40736 56176
rect 40972 55962 41000 56306
rect 41064 56273 41092 56494
rect 41340 56370 41368 56646
rect 41328 56364 41380 56370
rect 41328 56306 41380 56312
rect 41050 56264 41106 56273
rect 41050 56199 41106 56208
rect 41144 56160 41196 56166
rect 41144 56102 41196 56108
rect 41604 56160 41656 56166
rect 41604 56102 41656 56108
rect 40960 55956 41012 55962
rect 40960 55898 41012 55904
rect 40592 55888 40644 55894
rect 41156 55865 41184 56102
rect 40592 55830 40644 55836
rect 41142 55856 41198 55865
rect 40604 55078 40632 55830
rect 41142 55791 41198 55800
rect 41616 55758 41644 56102
rect 41708 55865 41736 59214
rect 41878 59200 41934 60000
rect 42338 59200 42394 60000
rect 42798 59200 42854 60000
rect 43258 59200 43314 60000
rect 43718 59200 43774 60000
rect 44178 59200 44234 60000
rect 44638 59200 44694 60000
rect 45098 59200 45154 60000
rect 45558 59200 45614 60000
rect 46018 59200 46074 60000
rect 46478 59200 46534 60000
rect 46584 59214 46888 59242
rect 41788 56840 41840 56846
rect 41788 56782 41840 56788
rect 41694 55856 41750 55865
rect 41800 55826 41828 56782
rect 41892 56409 41920 59200
rect 42156 56772 42208 56778
rect 42156 56714 42208 56720
rect 42064 56500 42116 56506
rect 42064 56442 42116 56448
rect 41878 56400 41934 56409
rect 41878 56335 41934 56344
rect 41694 55791 41750 55800
rect 41788 55820 41840 55826
rect 41788 55762 41840 55768
rect 41604 55752 41656 55758
rect 41604 55694 41656 55700
rect 41420 55616 41472 55622
rect 41420 55558 41472 55564
rect 40592 55072 40644 55078
rect 40592 55014 40644 55020
rect 40776 55072 40828 55078
rect 40776 55014 40828 55020
rect 40788 54670 40816 55014
rect 40500 54664 40552 54670
rect 40500 54606 40552 54612
rect 40776 54664 40828 54670
rect 40776 54606 40828 54612
rect 41328 54664 41380 54670
rect 41328 54606 41380 54612
rect 40408 54256 40460 54262
rect 40408 54198 40460 54204
rect 40316 54188 40368 54194
rect 40316 54130 40368 54136
rect 40040 54052 40092 54058
rect 40040 53994 40092 54000
rect 40420 53786 40448 54198
rect 40512 53990 40540 54606
rect 41340 54330 41368 54606
rect 41432 54602 41460 55558
rect 41420 54596 41472 54602
rect 41420 54538 41472 54544
rect 41328 54324 41380 54330
rect 41328 54266 41380 54272
rect 41432 54194 41460 54538
rect 41616 54262 41644 55694
rect 41800 55418 41828 55762
rect 41972 55616 42024 55622
rect 41972 55558 42024 55564
rect 41788 55412 41840 55418
rect 41788 55354 41840 55360
rect 41604 54256 41656 54262
rect 41604 54198 41656 54204
rect 41420 54188 41472 54194
rect 41420 54130 41472 54136
rect 41984 53990 42012 55558
rect 42076 54874 42104 56442
rect 42168 56370 42196 56714
rect 42352 56545 42380 59200
rect 42812 57974 42840 59200
rect 42812 57946 42932 57974
rect 42904 57390 42932 57946
rect 42892 57384 42944 57390
rect 42892 57326 42944 57332
rect 43076 57384 43128 57390
rect 43076 57326 43128 57332
rect 42708 56840 42760 56846
rect 42708 56782 42760 56788
rect 42338 56536 42394 56545
rect 42338 56471 42394 56480
rect 42156 56364 42208 56370
rect 42156 56306 42208 56312
rect 42720 56166 42748 56782
rect 42800 56228 42852 56234
rect 42800 56170 42852 56176
rect 42708 56160 42760 56166
rect 42708 56102 42760 56108
rect 42812 56001 42840 56170
rect 42798 55992 42854 56001
rect 42798 55927 42854 55936
rect 42248 55752 42300 55758
rect 42248 55694 42300 55700
rect 42524 55752 42576 55758
rect 42524 55694 42576 55700
rect 42260 55078 42288 55694
rect 42536 55418 42564 55694
rect 42616 55684 42668 55690
rect 42616 55626 42668 55632
rect 42524 55412 42576 55418
rect 42524 55354 42576 55360
rect 42536 55282 42564 55354
rect 42524 55276 42576 55282
rect 42524 55218 42576 55224
rect 42248 55072 42300 55078
rect 42248 55014 42300 55020
rect 42064 54868 42116 54874
rect 42064 54810 42116 54816
rect 42260 54330 42288 55014
rect 42536 54670 42564 55218
rect 42628 55214 42656 55626
rect 42616 55208 42668 55214
rect 42616 55150 42668 55156
rect 42524 54664 42576 54670
rect 42524 54606 42576 54612
rect 42904 54330 42932 57326
rect 42984 56296 43036 56302
rect 42984 56238 43036 56244
rect 42996 54670 43024 56238
rect 43088 55690 43116 57326
rect 43168 56704 43220 56710
rect 43168 56646 43220 56652
rect 43180 56370 43208 56646
rect 43168 56364 43220 56370
rect 43168 56306 43220 56312
rect 43076 55684 43128 55690
rect 43076 55626 43128 55632
rect 43088 55350 43116 55626
rect 43076 55344 43128 55350
rect 43076 55286 43128 55292
rect 42984 54664 43036 54670
rect 42984 54606 43036 54612
rect 43180 54602 43208 56306
rect 43272 54874 43300 59200
rect 43444 57928 43496 57934
rect 43444 57870 43496 57876
rect 43456 56846 43484 57870
rect 43444 56840 43496 56846
rect 43444 56782 43496 56788
rect 43732 56370 43760 59200
rect 43812 57588 43864 57594
rect 43812 57530 43864 57536
rect 43996 57588 44048 57594
rect 43996 57530 44048 57536
rect 43824 57390 43852 57530
rect 43812 57384 43864 57390
rect 43812 57326 43864 57332
rect 43824 56982 43852 57326
rect 43812 56976 43864 56982
rect 43812 56918 43864 56924
rect 43720 56364 43772 56370
rect 43720 56306 43772 56312
rect 43720 56228 43772 56234
rect 43720 56170 43772 56176
rect 43350 55856 43406 55865
rect 43350 55791 43352 55800
rect 43404 55791 43406 55800
rect 43352 55762 43404 55768
rect 43628 55752 43680 55758
rect 43628 55694 43680 55700
rect 43640 55622 43668 55694
rect 43732 55622 43760 56170
rect 43824 55758 43852 56918
rect 44008 56370 44036 57530
rect 44192 57338 44220 59200
rect 44548 57384 44600 57390
rect 44192 57310 44312 57338
rect 44548 57326 44600 57332
rect 44180 57248 44232 57254
rect 44180 57190 44232 57196
rect 44192 56914 44220 57190
rect 44180 56908 44232 56914
rect 44180 56850 44232 56856
rect 44088 56840 44140 56846
rect 44140 56788 44220 56794
rect 44088 56782 44220 56788
rect 44100 56766 44220 56782
rect 44088 56432 44140 56438
rect 44088 56374 44140 56380
rect 43996 56364 44048 56370
rect 43916 56324 43996 56352
rect 43812 55752 43864 55758
rect 43812 55694 43864 55700
rect 43628 55616 43680 55622
rect 43628 55558 43680 55564
rect 43720 55616 43772 55622
rect 43720 55558 43772 55564
rect 43260 54868 43312 54874
rect 43260 54810 43312 54816
rect 43168 54596 43220 54602
rect 43168 54538 43220 54544
rect 42248 54324 42300 54330
rect 42248 54266 42300 54272
rect 42892 54324 42944 54330
rect 42892 54266 42944 54272
rect 43732 54194 43760 55558
rect 43916 55282 43944 56324
rect 43996 56306 44048 56312
rect 44100 56234 44128 56374
rect 44192 56234 44220 56766
rect 44088 56228 44140 56234
rect 44088 56170 44140 56176
rect 44180 56228 44232 56234
rect 44180 56170 44232 56176
rect 43904 55276 43956 55282
rect 43904 55218 43956 55224
rect 44100 55214 44128 56170
rect 44192 55282 44220 56170
rect 44284 55350 44312 57310
rect 44364 56364 44416 56370
rect 44364 56306 44416 56312
rect 44376 55962 44404 56306
rect 44364 55956 44416 55962
rect 44364 55898 44416 55904
rect 44376 55418 44404 55898
rect 44560 55457 44588 57326
rect 44652 55962 44680 59200
rect 44824 57792 44876 57798
rect 44824 57734 44876 57740
rect 44732 57384 44784 57390
rect 44732 57326 44784 57332
rect 44744 56846 44772 57326
rect 44732 56840 44784 56846
rect 44732 56782 44784 56788
rect 44836 56370 44864 57734
rect 45008 57248 45060 57254
rect 45008 57190 45060 57196
rect 45020 56914 45048 57190
rect 45008 56908 45060 56914
rect 45008 56850 45060 56856
rect 45112 56370 45140 59200
rect 45572 57526 45600 59200
rect 45560 57520 45612 57526
rect 45560 57462 45612 57468
rect 45836 57520 45888 57526
rect 45836 57462 45888 57468
rect 45744 57248 45796 57254
rect 45744 57190 45796 57196
rect 45650 56944 45706 56953
rect 45650 56879 45706 56888
rect 45664 56846 45692 56879
rect 45652 56840 45704 56846
rect 45652 56782 45704 56788
rect 45468 56704 45520 56710
rect 45466 56672 45468 56681
rect 45520 56672 45522 56681
rect 45466 56607 45522 56616
rect 44824 56364 44876 56370
rect 44824 56306 44876 56312
rect 45100 56364 45152 56370
rect 45100 56306 45152 56312
rect 45560 56296 45612 56302
rect 45558 56264 45560 56273
rect 45612 56264 45614 56273
rect 45558 56199 45614 56208
rect 44824 56160 44876 56166
rect 44824 56102 44876 56108
rect 44640 55956 44692 55962
rect 44640 55898 44692 55904
rect 44836 55622 44864 56102
rect 44916 55888 44968 55894
rect 45100 55888 45152 55894
rect 44968 55848 45100 55876
rect 44916 55830 44968 55836
rect 45100 55830 45152 55836
rect 45560 55752 45612 55758
rect 45560 55694 45612 55700
rect 44824 55616 44876 55622
rect 44824 55558 44876 55564
rect 44546 55448 44602 55457
rect 44364 55412 44416 55418
rect 44546 55383 44602 55392
rect 44730 55448 44786 55457
rect 45572 55418 45600 55694
rect 45664 55418 45692 56782
rect 45756 56438 45784 57190
rect 45744 56432 45796 56438
rect 45744 56374 45796 56380
rect 45848 55962 45876 57462
rect 46032 57050 46060 59200
rect 46492 59106 46520 59200
rect 46584 59106 46612 59214
rect 46492 59078 46612 59106
rect 46860 57066 46888 59214
rect 46938 59200 46994 60000
rect 47398 59200 47454 60000
rect 47858 59200 47914 60000
rect 48318 59200 48374 60000
rect 48778 59200 48834 60000
rect 49238 59200 49294 60000
rect 49344 59214 49648 59242
rect 46952 57458 46980 59200
rect 46940 57452 46992 57458
rect 46992 57412 47072 57440
rect 46940 57394 46992 57400
rect 46020 57044 46072 57050
rect 46860 57038 46980 57066
rect 46020 56986 46072 56992
rect 46952 56982 46980 57038
rect 46940 56976 46992 56982
rect 46940 56918 46992 56924
rect 46112 56840 46164 56846
rect 46112 56782 46164 56788
rect 46940 56840 46992 56846
rect 46940 56782 46992 56788
rect 46124 56409 46152 56782
rect 46952 56545 46980 56782
rect 46938 56536 46994 56545
rect 46938 56471 46994 56480
rect 46110 56400 46166 56409
rect 46110 56335 46166 56344
rect 47044 55962 47072 57412
rect 47216 57384 47268 57390
rect 47216 57326 47268 57332
rect 47228 56166 47256 57326
rect 47412 56370 47440 59200
rect 47872 56370 47900 59200
rect 48332 57458 48360 59200
rect 48320 57452 48372 57458
rect 48320 57394 48372 57400
rect 48332 56506 48360 57394
rect 48792 57050 48820 59200
rect 49252 59106 49280 59200
rect 49344 59106 49372 59214
rect 49252 59078 49372 59106
rect 49620 57236 49648 59214
rect 49698 59200 49754 60000
rect 50158 59200 50214 60000
rect 50618 59200 50674 60000
rect 51078 59200 51134 60000
rect 51538 59200 51594 60000
rect 51998 59200 52054 60000
rect 52104 59214 52408 59242
rect 49712 57458 49740 59200
rect 49700 57452 49752 57458
rect 49752 57412 49832 57440
rect 49700 57394 49752 57400
rect 49620 57208 49740 57236
rect 49712 57050 49740 57208
rect 48780 57044 48832 57050
rect 48780 56986 48832 56992
rect 49700 57044 49752 57050
rect 49700 56986 49752 56992
rect 49804 56506 49832 57412
rect 50068 57316 50120 57322
rect 50068 57258 50120 57264
rect 48320 56500 48372 56506
rect 48320 56442 48372 56448
rect 49792 56500 49844 56506
rect 49792 56442 49844 56448
rect 47400 56364 47452 56370
rect 47400 56306 47452 56312
rect 47860 56364 47912 56370
rect 47860 56306 47912 56312
rect 47216 56160 47268 56166
rect 47216 56102 47268 56108
rect 45836 55956 45888 55962
rect 45836 55898 45888 55904
rect 47032 55956 47084 55962
rect 47032 55898 47084 55904
rect 50080 55826 50108 57258
rect 50172 57050 50200 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 50632 57050 50660 59200
rect 51092 57458 51120 59200
rect 51264 57860 51316 57866
rect 51264 57802 51316 57808
rect 51276 57594 51304 57802
rect 51264 57588 51316 57594
rect 51264 57530 51316 57536
rect 51080 57452 51132 57458
rect 51080 57394 51132 57400
rect 51080 57248 51132 57254
rect 51080 57190 51132 57196
rect 50160 57044 50212 57050
rect 50160 56986 50212 56992
rect 50620 57044 50672 57050
rect 50620 56986 50672 56992
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 51092 55894 51120 57190
rect 51552 57050 51580 59200
rect 52012 59106 52040 59200
rect 52104 59106 52132 59214
rect 52012 59078 52132 59106
rect 51632 57452 51684 57458
rect 52380 57440 52408 59214
rect 52458 59200 52514 60000
rect 52918 59200 52974 60000
rect 53378 59200 53434 60000
rect 53838 59200 53894 60000
rect 54298 59200 54354 60000
rect 54758 59200 54814 60000
rect 55218 59200 55274 60000
rect 55678 59200 55734 60000
rect 56138 59200 56194 60000
rect 52472 57594 52500 59200
rect 52460 57588 52512 57594
rect 52460 57530 52512 57536
rect 52552 57520 52604 57526
rect 52552 57462 52604 57468
rect 52380 57412 52500 57440
rect 51632 57394 51684 57400
rect 51540 57044 51592 57050
rect 51540 56986 51592 56992
rect 51644 56506 51672 57394
rect 52472 57050 52500 57412
rect 52460 57044 52512 57050
rect 52460 56986 52512 56992
rect 52564 56506 52592 57462
rect 52932 57050 52960 59200
rect 53392 57050 53420 59200
rect 53852 57458 53880 59200
rect 53840 57452 53892 57458
rect 53840 57394 53892 57400
rect 52920 57044 52972 57050
rect 52920 56986 52972 56992
rect 53380 57044 53432 57050
rect 53380 56986 53432 56992
rect 53852 56506 53880 57394
rect 54116 57248 54168 57254
rect 54116 57190 54168 57196
rect 54128 56982 54156 57190
rect 54312 57050 54340 59200
rect 54300 57044 54352 57050
rect 54300 56986 54352 56992
rect 54116 56976 54168 56982
rect 54116 56918 54168 56924
rect 54772 56914 54800 59200
rect 55232 57458 55260 59200
rect 55692 57458 55720 59200
rect 55220 57452 55272 57458
rect 55220 57394 55272 57400
rect 55680 57452 55732 57458
rect 55680 57394 55732 57400
rect 54760 56908 54812 56914
rect 54760 56850 54812 56856
rect 55232 56506 55260 57394
rect 56152 57050 56180 59200
rect 56140 57044 56192 57050
rect 56140 56986 56192 56992
rect 51632 56500 51684 56506
rect 51632 56442 51684 56448
rect 52552 56500 52604 56506
rect 52552 56442 52604 56448
rect 53840 56500 53892 56506
rect 53840 56442 53892 56448
rect 55220 56500 55272 56506
rect 55220 56442 55272 56448
rect 51080 55888 51132 55894
rect 51080 55830 51132 55836
rect 50068 55820 50120 55826
rect 50068 55762 50120 55768
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 44730 55383 44732 55392
rect 44364 55354 44416 55360
rect 44784 55383 44786 55392
rect 45560 55412 45612 55418
rect 44732 55354 44784 55360
rect 45560 55354 45612 55360
rect 45652 55412 45704 55418
rect 45652 55354 45704 55360
rect 44272 55344 44324 55350
rect 44272 55286 44324 55292
rect 44180 55276 44232 55282
rect 44180 55218 44232 55224
rect 44088 55208 44140 55214
rect 44088 55150 44140 55156
rect 44284 54874 44312 55286
rect 44272 54868 44324 54874
rect 44272 54810 44324 54816
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 43720 54188 43772 54194
rect 43720 54130 43772 54136
rect 40500 53984 40552 53990
rect 40500 53926 40552 53932
rect 41972 53984 42024 53990
rect 41972 53926 42024 53932
rect 40408 53780 40460 53786
rect 40408 53722 40460 53728
rect 39856 53712 39908 53718
rect 39856 53654 39908 53660
rect 36452 53644 36504 53650
rect 36452 53586 36504 53592
rect 40420 53242 40448 53722
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 36084 53236 36136 53242
rect 36084 53178 36136 53184
rect 40408 53236 40460 53242
rect 40408 53178 40460 53184
rect 35992 52692 36044 52698
rect 35992 52634 36044 52640
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 34716 45526 34836 45554
rect 34716 12434 34744 45526
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34624 12406 34744 12434
rect 27712 8084 27764 8090
rect 27712 8026 27764 8032
rect 30840 8084 30892 8090
rect 30840 8026 30892 8032
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 26240 7404 26292 7410
rect 26240 7346 26292 7352
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 26252 6798 26280 7346
rect 27436 7200 27488 7206
rect 27436 7142 27488 7148
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26608 6792 26660 6798
rect 26608 6734 26660 6740
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 25148 6458 25176 6598
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 24308 5704 24360 5710
rect 24308 5646 24360 5652
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 7668 800 7696 2382
rect 8220 800 8248 2382
rect 8588 800 8616 2790
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 8956 800 8984 2382
rect 9324 800 9352 2790
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9692 800 9720 2382
rect 9968 800 9996 2790
rect 10244 800 10272 3470
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 10520 800 10548 2518
rect 10796 800 10824 2790
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11072 800 11100 2382
rect 11348 800 11376 2790
rect 11624 800 11652 2790
rect 11888 2576 11940 2582
rect 11888 2518 11940 2524
rect 11900 800 11928 2518
rect 12176 800 12204 3470
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12452 800 12480 2382
rect 12728 800 12756 2790
rect 13004 800 13032 3470
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 13280 800 13308 2518
rect 13556 800 13584 2790
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 13832 800 13860 2382
rect 14108 800 14136 3470
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 14384 800 14412 2790
rect 14648 2576 14700 2582
rect 14648 2518 14700 2524
rect 14660 800 14688 2518
rect 14936 800 14964 3470
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15212 800 15240 2790
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15488 800 15516 2382
rect 15764 800 15792 3470
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 16040 800 16068 2790
rect 16316 800 16344 2790
rect 16592 800 16620 3470
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 16868 800 16896 2450
rect 17144 800 17172 3878
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17328 800 17356 2790
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17604 800 17632 2518
rect 17880 800 17908 3470
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18156 800 18184 2586
rect 18432 800 18460 3878
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 18708 800 18736 3470
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 18984 800 19012 2926
rect 19260 800 19288 3470
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 19352 1306 19380 2450
rect 19444 1442 19472 2858
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 2106 20024 2382
rect 19984 2100 20036 2106
rect 19984 2042 20036 2048
rect 19444 1414 19840 1442
rect 19352 1278 19564 1306
rect 19536 800 19564 1278
rect 19812 800 19840 1414
rect 20088 800 20116 3878
rect 20364 800 20392 3878
rect 20732 2802 20760 4558
rect 21732 3664 21784 3670
rect 21732 3606 21784 3612
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 20640 2774 20760 2802
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 20640 800 20668 2774
rect 20916 800 20944 2790
rect 21192 800 21220 3538
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 21376 2038 21404 2382
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 21364 2032 21416 2038
rect 21364 1974 21416 1980
rect 21468 800 21496 2314
rect 21744 800 21772 3606
rect 22020 800 22048 4558
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22100 4004 22152 4010
rect 22100 3946 22152 3952
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 22112 3738 22140 3946
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 22112 3058 22140 3334
rect 22204 3194 22232 3946
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 22296 800 22324 4014
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22480 3602 22508 3878
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 22376 3528 22428 3534
rect 22376 3470 22428 3476
rect 22388 3058 22416 3470
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 22572 800 22600 4966
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22664 3602 22692 4422
rect 22652 3596 22704 3602
rect 22652 3538 22704 3544
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 22756 2774 22784 2858
rect 22756 2746 22876 2774
rect 22744 2644 22796 2650
rect 22744 2586 22796 2592
rect 22756 2310 22784 2586
rect 22744 2304 22796 2310
rect 22744 2246 22796 2252
rect 22848 800 22876 2746
rect 23112 2576 23164 2582
rect 23112 2518 23164 2524
rect 23124 800 23152 2518
rect 23400 800 23428 5646
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 23940 4752 23992 4758
rect 23940 4694 23992 4700
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23492 4146 23520 4558
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23492 3398 23520 4082
rect 23848 4072 23900 4078
rect 23848 4014 23900 4020
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23492 2446 23520 3334
rect 23860 2650 23888 4014
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23664 2100 23716 2106
rect 23664 2042 23716 2048
rect 23676 800 23704 2042
rect 23952 800 23980 4694
rect 24044 3126 24072 5510
rect 24320 5234 24348 5646
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24320 4622 24348 5170
rect 24872 5166 24900 6190
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 24860 5160 24912 5166
rect 24860 5102 24912 5108
rect 24308 4616 24360 4622
rect 24308 4558 24360 4564
rect 24964 3738 24992 5646
rect 25240 4690 25268 6734
rect 25688 6316 25740 6322
rect 25688 6258 25740 6264
rect 25412 6112 25464 6118
rect 25412 6054 25464 6060
rect 25424 4690 25452 6054
rect 25504 5636 25556 5642
rect 25504 5578 25556 5584
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 25228 4684 25280 4690
rect 25228 4626 25280 4632
rect 25412 4684 25464 4690
rect 25412 4626 25464 4632
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 25056 3602 25084 4626
rect 25320 4140 25372 4146
rect 25320 4082 25372 4088
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 25148 3738 25176 3878
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 25044 3596 25096 3602
rect 25044 3538 25096 3544
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24032 3120 24084 3126
rect 24032 3062 24084 3068
rect 24228 800 24256 3402
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 24504 800 24532 3130
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24768 2372 24820 2378
rect 24768 2314 24820 2320
rect 24780 800 24808 2314
rect 24872 1426 24900 2450
rect 24860 1420 24912 1426
rect 24860 1362 24912 1368
rect 25056 800 25084 2926
rect 25332 2650 25360 4082
rect 25412 3460 25464 3466
rect 25412 3402 25464 3408
rect 25320 2644 25372 2650
rect 25320 2586 25372 2592
rect 25424 2582 25452 3402
rect 25516 2922 25544 5578
rect 25700 5234 25728 6258
rect 26252 5386 26280 6734
rect 26160 5358 26280 5386
rect 26160 5302 26188 5358
rect 26148 5296 26200 5302
rect 26148 5238 26200 5244
rect 26620 5234 26648 6734
rect 26792 6656 26844 6662
rect 26792 6598 26844 6604
rect 26804 6390 26832 6598
rect 26792 6384 26844 6390
rect 26792 6326 26844 6332
rect 26700 5772 26752 5778
rect 26700 5714 26752 5720
rect 25688 5228 25740 5234
rect 25688 5170 25740 5176
rect 26608 5228 26660 5234
rect 26608 5170 26660 5176
rect 26240 4684 26292 4690
rect 26240 4626 26292 4632
rect 26148 4480 26200 4486
rect 26148 4422 26200 4428
rect 26160 3670 26188 4422
rect 26148 3664 26200 3670
rect 26148 3606 26200 3612
rect 25504 2916 25556 2922
rect 25504 2858 25556 2864
rect 26252 2774 26280 4626
rect 26516 4004 26568 4010
rect 26516 3946 26568 3952
rect 26424 3392 26476 3398
rect 26424 3334 26476 3340
rect 26160 2746 26280 2774
rect 25412 2576 25464 2582
rect 25412 2518 25464 2524
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25320 2032 25372 2038
rect 25320 1974 25372 1980
rect 25332 800 25360 1974
rect 25596 1420 25648 1426
rect 25596 1362 25648 1368
rect 25608 800 25636 1362
rect 25884 800 25912 2246
rect 26160 800 26188 2746
rect 26436 800 26464 3334
rect 26528 2514 26556 3946
rect 26608 2984 26660 2990
rect 26608 2926 26660 2932
rect 26620 2650 26648 2926
rect 26608 2644 26660 2650
rect 26608 2586 26660 2592
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 26712 800 26740 5714
rect 27448 5302 27476 7142
rect 27620 6792 27672 6798
rect 27620 6734 27672 6740
rect 27528 6248 27580 6254
rect 27528 6190 27580 6196
rect 27436 5296 27488 5302
rect 27436 5238 27488 5244
rect 26976 3936 27028 3942
rect 26976 3878 27028 3884
rect 26792 2984 26844 2990
rect 26792 2926 26844 2932
rect 26804 2582 26832 2926
rect 26792 2576 26844 2582
rect 26792 2518 26844 2524
rect 26988 800 27016 3878
rect 27252 3120 27304 3126
rect 27252 3062 27304 3068
rect 27264 800 27292 3062
rect 27540 800 27568 6190
rect 27632 4690 27660 6734
rect 27724 6458 27752 8026
rect 29644 7880 29696 7886
rect 29644 7822 29696 7828
rect 29552 7744 29604 7750
rect 29552 7686 29604 7692
rect 27988 7200 28040 7206
rect 27988 7142 28040 7148
rect 29460 7200 29512 7206
rect 29460 7142 29512 7148
rect 27712 6452 27764 6458
rect 27712 6394 27764 6400
rect 27896 5704 27948 5710
rect 27896 5646 27948 5652
rect 27712 5160 27764 5166
rect 27712 5102 27764 5108
rect 27620 4684 27672 4690
rect 27620 4626 27672 4632
rect 27724 2632 27752 5102
rect 27804 5024 27856 5030
rect 27804 4966 27856 4972
rect 27816 4690 27844 4966
rect 27804 4684 27856 4690
rect 27804 4626 27856 4632
rect 27908 2854 27936 5646
rect 28000 3602 28028 7142
rect 29000 6792 29052 6798
rect 29000 6734 29052 6740
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29368 6792 29420 6798
rect 29368 6734 29420 6740
rect 28632 5772 28684 5778
rect 28632 5714 28684 5720
rect 28080 5636 28132 5642
rect 28080 5578 28132 5584
rect 28092 3738 28120 5578
rect 28172 4684 28224 4690
rect 28172 4626 28224 4632
rect 28080 3732 28132 3738
rect 28080 3674 28132 3680
rect 27988 3596 28040 3602
rect 27988 3538 28040 3544
rect 27896 2848 27948 2854
rect 27896 2790 27948 2796
rect 27724 2604 27844 2632
rect 27816 800 27844 2604
rect 28184 2292 28212 4626
rect 28356 3596 28408 3602
rect 28356 3538 28408 3544
rect 28092 2264 28212 2292
rect 28092 800 28120 2264
rect 28368 800 28396 3538
rect 28540 2984 28592 2990
rect 28540 2926 28592 2932
rect 28552 2650 28580 2926
rect 28540 2644 28592 2650
rect 28540 2586 28592 2592
rect 28644 800 28672 5714
rect 29012 4146 29040 6734
rect 29288 6322 29316 6734
rect 29276 6316 29328 6322
rect 29276 6258 29328 6264
rect 29380 5234 29408 6734
rect 29472 6390 29500 7142
rect 29460 6384 29512 6390
rect 29460 6326 29512 6332
rect 29368 5228 29420 5234
rect 29368 5170 29420 5176
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 29564 4078 29592 7686
rect 29656 7410 29684 7822
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29656 6730 29684 7346
rect 30196 7200 30248 7206
rect 30196 7142 30248 7148
rect 29644 6724 29696 6730
rect 29644 6666 29696 6672
rect 29552 4072 29604 4078
rect 29552 4014 29604 4020
rect 29184 4004 29236 4010
rect 29184 3946 29236 3952
rect 28908 3460 28960 3466
rect 28908 3402 28960 3408
rect 28920 800 28948 3402
rect 29196 800 29224 3946
rect 29552 2984 29604 2990
rect 29552 2926 29604 2932
rect 29460 2916 29512 2922
rect 29460 2858 29512 2864
rect 29472 800 29500 2858
rect 29564 2582 29592 2926
rect 29552 2576 29604 2582
rect 29552 2518 29604 2524
rect 29656 2446 29684 6666
rect 30012 6248 30064 6254
rect 30012 6190 30064 6196
rect 29736 4072 29788 4078
rect 29736 4014 29788 4020
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 29748 800 29776 4014
rect 30024 800 30052 6190
rect 30208 5302 30236 7142
rect 30852 6798 30880 8026
rect 32036 7404 32088 7410
rect 32036 7346 32088 7352
rect 32956 7404 33008 7410
rect 32956 7346 33008 7352
rect 30932 7200 30984 7206
rect 30932 7142 30984 7148
rect 30840 6792 30892 6798
rect 30840 6734 30892 6740
rect 30852 6322 30880 6734
rect 30840 6316 30892 6322
rect 30840 6258 30892 6264
rect 30944 5778 30972 7142
rect 32048 6866 32076 7346
rect 32312 7200 32364 7206
rect 32312 7142 32364 7148
rect 32036 6860 32088 6866
rect 32036 6802 32088 6808
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 31772 5846 31800 6734
rect 32036 6724 32088 6730
rect 32036 6666 32088 6672
rect 32048 6390 32076 6666
rect 32036 6384 32088 6390
rect 32036 6326 32088 6332
rect 32128 6112 32180 6118
rect 32128 6054 32180 6060
rect 31760 5840 31812 5846
rect 31760 5782 31812 5788
rect 30932 5772 30984 5778
rect 30932 5714 30984 5720
rect 31668 5772 31720 5778
rect 31668 5714 31720 5720
rect 30196 5296 30248 5302
rect 30196 5238 30248 5244
rect 30380 5160 30432 5166
rect 30380 5102 30432 5108
rect 30392 4706 30420 5102
rect 30300 4678 30420 4706
rect 30748 4684 30800 4690
rect 30300 800 30328 4678
rect 30748 4626 30800 4632
rect 30380 4616 30432 4622
rect 30432 4576 30512 4604
rect 30380 4558 30432 4564
rect 30380 3460 30432 3466
rect 30380 3402 30432 3408
rect 30392 2650 30420 3402
rect 30380 2644 30432 2650
rect 30380 2586 30432 2592
rect 30484 2514 30512 4576
rect 30656 4548 30708 4554
rect 30656 4490 30708 4496
rect 30564 3528 30616 3534
rect 30564 3470 30616 3476
rect 30576 2650 30604 3470
rect 30564 2644 30616 2650
rect 30564 2586 30616 2592
rect 30472 2508 30524 2514
rect 30472 2450 30524 2456
rect 30668 2378 30696 4490
rect 30656 2372 30708 2378
rect 30656 2314 30708 2320
rect 30760 2258 30788 4626
rect 30840 3596 30892 3602
rect 30840 3538 30892 3544
rect 30576 2230 30788 2258
rect 30576 800 30604 2230
rect 30852 800 30880 3538
rect 31116 2984 31168 2990
rect 31116 2926 31168 2932
rect 31128 800 31156 2926
rect 31392 2848 31444 2854
rect 31392 2790 31444 2796
rect 31404 800 31432 2790
rect 31680 800 31708 5714
rect 31760 5160 31812 5166
rect 31760 5102 31812 5108
rect 31772 2854 31800 5102
rect 32140 4146 32168 6054
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 32324 4078 32352 7142
rect 32968 6322 32996 7346
rect 33232 7200 33284 7206
rect 33232 7142 33284 7148
rect 33140 6792 33192 6798
rect 33140 6734 33192 6740
rect 32956 6316 33008 6322
rect 32956 6258 33008 6264
rect 32312 4072 32364 4078
rect 32312 4014 32364 4020
rect 32772 4072 32824 4078
rect 32772 4014 32824 4020
rect 32220 3596 32272 3602
rect 32220 3538 32272 3544
rect 31944 2984 31996 2990
rect 31944 2926 31996 2932
rect 31760 2848 31812 2854
rect 31760 2790 31812 2796
rect 31956 800 31984 2926
rect 32232 800 32260 3538
rect 32496 2916 32548 2922
rect 32496 2858 32548 2864
rect 32508 800 32536 2858
rect 32784 800 32812 4014
rect 32968 2446 32996 6258
rect 33152 4690 33180 6734
rect 33244 4758 33272 7142
rect 33968 6792 34020 6798
rect 33968 6734 34020 6740
rect 33416 6656 33468 6662
rect 33416 6598 33468 6604
rect 33324 5772 33376 5778
rect 33324 5714 33376 5720
rect 33232 4752 33284 4758
rect 33232 4694 33284 4700
rect 33140 4684 33192 4690
rect 33140 4626 33192 4632
rect 33140 3528 33192 3534
rect 33140 3470 33192 3476
rect 33048 3188 33100 3194
rect 33048 3130 33100 3136
rect 32956 2440 33008 2446
rect 32956 2382 33008 2388
rect 33060 800 33088 3130
rect 33152 2650 33180 3470
rect 33140 2644 33192 2650
rect 33140 2586 33192 2592
rect 33336 800 33364 5714
rect 33428 5302 33456 6598
rect 33600 6180 33652 6186
rect 33600 6122 33652 6128
rect 33416 5296 33468 5302
rect 33416 5238 33468 5244
rect 33612 5234 33640 6122
rect 33980 5846 34008 6734
rect 33968 5840 34020 5846
rect 33968 5782 34020 5788
rect 33600 5228 33652 5234
rect 33600 5170 33652 5176
rect 34520 5160 34572 5166
rect 34520 5102 34572 5108
rect 33600 4684 33652 4690
rect 33600 4626 33652 4632
rect 33612 3194 33640 4626
rect 34060 4072 34112 4078
rect 34532 4026 34560 5102
rect 34060 4014 34112 4020
rect 33692 3596 33744 3602
rect 33692 3538 33744 3544
rect 33600 3188 33652 3194
rect 33600 3130 33652 3136
rect 33416 2984 33468 2990
rect 33416 2926 33468 2932
rect 33600 2984 33652 2990
rect 33600 2926 33652 2932
rect 33428 2650 33456 2926
rect 33416 2644 33468 2650
rect 33416 2586 33468 2592
rect 33612 2582 33640 2926
rect 33600 2576 33652 2582
rect 33600 2518 33652 2524
rect 33704 1850 33732 3538
rect 33876 3460 33928 3466
rect 33876 3402 33928 3408
rect 33888 2650 33916 3402
rect 33876 2644 33928 2650
rect 33876 2586 33928 2592
rect 34072 2122 34100 4014
rect 34440 3998 34560 4026
rect 34152 3120 34204 3126
rect 34152 3062 34204 3068
rect 33612 1822 33732 1850
rect 33888 2094 34100 2122
rect 33612 800 33640 1822
rect 33888 800 33916 2094
rect 34164 800 34192 3062
rect 34440 800 34468 3998
rect 34520 2984 34572 2990
rect 34520 2926 34572 2932
rect 34532 2650 34560 2926
rect 34520 2644 34572 2650
rect 34520 2586 34572 2592
rect 34624 2530 34652 12406
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 34796 6112 34848 6118
rect 34796 6054 34848 6060
rect 34808 5778 34836 6054
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34796 5772 34848 5778
rect 34796 5714 34848 5720
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 37924 5296 37976 5302
rect 37924 5238 37976 5244
rect 37188 5160 37240 5166
rect 37188 5102 37240 5108
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 37200 4826 37228 5102
rect 37188 4820 37240 4826
rect 37188 4762 37240 4768
rect 36360 4616 36412 4622
rect 36360 4558 36412 4564
rect 36728 4616 36780 4622
rect 36728 4558 36780 4564
rect 37832 4616 37884 4622
rect 37832 4558 37884 4564
rect 36176 4480 36228 4486
rect 36176 4422 36228 4428
rect 36188 4214 36216 4422
rect 36176 4208 36228 4214
rect 36176 4150 36228 4156
rect 36372 4146 36400 4558
rect 36360 4140 36412 4146
rect 36360 4082 36412 4088
rect 35808 4072 35860 4078
rect 35808 4014 35860 4020
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35532 3392 35584 3398
rect 35532 3334 35584 3340
rect 35348 3188 35400 3194
rect 35348 3130 35400 3136
rect 34704 2984 34756 2990
rect 34704 2926 34756 2932
rect 34716 2650 34744 2926
rect 34796 2848 34848 2854
rect 34796 2790 34848 2796
rect 34704 2644 34756 2650
rect 34704 2586 34756 2592
rect 34624 2502 34744 2530
rect 34716 800 34744 2502
rect 34808 1986 34836 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34808 1958 35020 1986
rect 34992 800 35020 1958
rect 35360 1170 35388 3130
rect 35268 1142 35388 1170
rect 35268 800 35296 1142
rect 35544 800 35572 3334
rect 35820 800 35848 4014
rect 36176 3664 36228 3670
rect 36176 3606 36228 3612
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 35912 2582 35940 3470
rect 36084 3460 36136 3466
rect 36084 3402 36136 3408
rect 36096 2650 36124 3402
rect 36084 2644 36136 2650
rect 36084 2586 36136 2592
rect 35900 2576 35952 2582
rect 35900 2518 35952 2524
rect 36188 1850 36216 3606
rect 36636 3460 36688 3466
rect 36636 3402 36688 3408
rect 36360 3120 36412 3126
rect 36360 3062 36412 3068
rect 36096 1822 36216 1850
rect 36096 800 36124 1822
rect 36372 800 36400 3062
rect 36648 800 36676 3402
rect 36740 2446 36768 4558
rect 37556 4004 37608 4010
rect 37556 3946 37608 3952
rect 37280 3936 37332 3942
rect 37280 3878 37332 3884
rect 36912 3732 36964 3738
rect 36912 3674 36964 3680
rect 36728 2440 36780 2446
rect 36728 2382 36780 2388
rect 36924 800 36952 3674
rect 37292 3058 37320 3878
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 37464 2984 37516 2990
rect 37464 2926 37516 2932
rect 37476 2650 37504 2926
rect 37464 2644 37516 2650
rect 37464 2586 37516 2592
rect 37188 2508 37240 2514
rect 37188 2450 37240 2456
rect 37200 800 37228 2450
rect 37568 1986 37596 3946
rect 37844 3738 37872 4558
rect 37832 3732 37884 3738
rect 37832 3674 37884 3680
rect 37936 2650 37964 5238
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 39120 4072 39172 4078
rect 39120 4014 39172 4020
rect 38292 3936 38344 3942
rect 38292 3878 38344 3884
rect 38016 2916 38068 2922
rect 38016 2858 38068 2864
rect 37924 2644 37976 2650
rect 37924 2586 37976 2592
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 37476 1958 37596 1986
rect 37476 800 37504 1958
rect 37752 800 37780 2314
rect 38028 800 38056 2858
rect 38304 800 38332 3878
rect 38568 3596 38620 3602
rect 38568 3538 38620 3544
rect 38580 800 38608 3538
rect 38844 3460 38896 3466
rect 38844 3402 38896 3408
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 38672 2650 38700 2790
rect 38660 2644 38712 2650
rect 38660 2586 38712 2592
rect 38856 800 38884 3402
rect 39132 800 39160 4014
rect 39948 4004 40000 4010
rect 39948 3946 40000 3952
rect 39304 3188 39356 3194
rect 39304 3130 39356 3136
rect 39316 2650 39344 3130
rect 39672 3052 39724 3058
rect 39672 2994 39724 3000
rect 39304 2644 39356 2650
rect 39304 2586 39356 2592
rect 39396 2576 39448 2582
rect 39396 2518 39448 2524
rect 39408 800 39436 2518
rect 39684 800 39712 2994
rect 39960 800 39988 3946
rect 40500 3664 40552 3670
rect 40500 3606 40552 3612
rect 42708 3664 42760 3670
rect 42708 3606 42760 3612
rect 40040 3392 40092 3398
rect 40040 3334 40092 3340
rect 40052 2650 40080 3334
rect 40224 2984 40276 2990
rect 40224 2926 40276 2932
rect 40040 2644 40092 2650
rect 40040 2586 40092 2592
rect 40236 800 40264 2926
rect 40512 800 40540 3606
rect 41328 3596 41380 3602
rect 41328 3538 41380 3544
rect 41052 2916 41104 2922
rect 41052 2858 41104 2864
rect 40776 2372 40828 2378
rect 40776 2314 40828 2320
rect 40788 800 40816 2314
rect 41064 800 41092 2858
rect 41340 800 41368 3538
rect 41880 3460 41932 3466
rect 41880 3402 41932 3408
rect 41604 2508 41656 2514
rect 41604 2450 41656 2456
rect 41616 800 41644 2450
rect 41892 800 41920 3402
rect 42156 2984 42208 2990
rect 42156 2926 42208 2932
rect 42168 800 42196 2926
rect 42432 2576 42484 2582
rect 42432 2518 42484 2524
rect 42444 800 42472 2518
rect 42720 800 42748 3606
rect 43536 3528 43588 3534
rect 43536 3470 43588 3476
rect 44916 3528 44968 3534
rect 44916 3470 44968 3476
rect 46296 3528 46348 3534
rect 46296 3470 46348 3476
rect 47676 3528 47728 3534
rect 47676 3470 47728 3476
rect 49056 3528 49108 3534
rect 49056 3470 49108 3476
rect 50620 3528 50672 3534
rect 50620 3470 50672 3476
rect 51816 3528 51868 3534
rect 51816 3470 51868 3476
rect 43260 2916 43312 2922
rect 43260 2858 43312 2864
rect 42984 2440 43036 2446
rect 42984 2382 43036 2388
rect 42996 800 43024 2382
rect 43272 800 43300 2858
rect 43548 800 43576 3470
rect 44640 2984 44692 2990
rect 44640 2926 44692 2932
rect 43812 2848 43864 2854
rect 43812 2790 43864 2796
rect 43824 800 43852 2790
rect 44088 2508 44140 2514
rect 44088 2450 44140 2456
rect 44100 800 44128 2450
rect 44364 2372 44416 2378
rect 44364 2314 44416 2320
rect 44376 800 44404 2314
rect 44652 800 44680 2926
rect 44928 800 44956 3470
rect 45468 2916 45520 2922
rect 45468 2858 45520 2864
rect 45192 2576 45244 2582
rect 45192 2518 45244 2524
rect 45204 800 45232 2518
rect 45480 800 45508 2858
rect 46020 2848 46072 2854
rect 46020 2790 46072 2796
rect 45744 2372 45796 2378
rect 45744 2314 45796 2320
rect 45756 800 45784 2314
rect 46032 800 46060 2790
rect 46308 800 46336 3470
rect 46572 2916 46624 2922
rect 46572 2858 46624 2864
rect 46584 800 46612 2858
rect 47400 2848 47452 2854
rect 47400 2790 47452 2796
rect 47124 2644 47176 2650
rect 47124 2586 47176 2592
rect 46848 2508 46900 2514
rect 46848 2450 46900 2456
rect 46860 800 46888 2450
rect 47136 800 47164 2586
rect 47412 800 47440 2790
rect 47688 800 47716 3470
rect 48228 2916 48280 2922
rect 48228 2858 48280 2864
rect 47952 2576 48004 2582
rect 47952 2518 48004 2524
rect 47964 800 47992 2518
rect 48240 800 48268 2858
rect 48780 2848 48832 2854
rect 48780 2790 48832 2796
rect 48504 2440 48556 2446
rect 48504 2382 48556 2388
rect 48516 800 48544 2382
rect 48792 800 48820 2790
rect 49068 800 49096 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 49332 2916 49384 2922
rect 49332 2858 49384 2864
rect 49344 800 49372 2858
rect 50160 2848 50212 2854
rect 50160 2790 50212 2796
rect 49884 2644 49936 2650
rect 49884 2586 49936 2592
rect 49608 2508 49660 2514
rect 49608 2450 49660 2456
rect 49620 800 49648 2450
rect 49896 800 49924 2586
rect 50172 800 50200 2790
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50632 1850 50660 3470
rect 50988 2916 51040 2922
rect 50988 2858 51040 2864
rect 50712 2372 50764 2378
rect 50712 2314 50764 2320
rect 50448 1822 50660 1850
rect 50448 800 50476 1822
rect 50724 800 50752 2314
rect 51000 800 51028 2858
rect 51540 2848 51592 2854
rect 51540 2790 51592 2796
rect 51264 2576 51316 2582
rect 51264 2518 51316 2524
rect 51276 800 51304 2518
rect 51552 800 51580 2790
rect 51828 800 51856 3470
rect 52092 2916 52144 2922
rect 52092 2858 52144 2864
rect 52104 800 52132 2858
rect 52368 2508 52420 2514
rect 52368 2450 52420 2456
rect 52380 800 52408 2450
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
<< via2 >>
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 6366 57452 6422 57488
rect 6366 57432 6368 57452
rect 6368 57432 6420 57452
rect 6420 57432 6422 57452
rect 11886 57296 11942 57352
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 20718 56888 20774 56944
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 25502 55800 25558 55856
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 27526 57704 27582 57760
rect 26882 56208 26938 56264
rect 27434 56888 27490 56944
rect 27526 56772 27582 56808
rect 27526 56752 27528 56772
rect 27528 56752 27580 56772
rect 27580 56752 27582 56772
rect 27710 57296 27766 57352
rect 27710 56616 27766 56672
rect 27986 57432 28042 57488
rect 28170 57704 28226 57760
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 29366 56364 29422 56400
rect 29366 56344 29368 56364
rect 29368 56344 29420 56364
rect 29420 56344 29422 56364
rect 29826 56616 29882 56672
rect 29826 56480 29882 56536
rect 29826 55392 29882 55448
rect 30010 56752 30066 56808
rect 32954 55392 33010 55448
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 36082 56480 36138 56536
rect 37370 56344 37426 56400
rect 37002 55936 37058 55992
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 37830 55936 37886 55992
rect 38014 55392 38070 55448
rect 40038 56888 40094 56944
rect 40590 56652 40592 56672
rect 40592 56652 40644 56672
rect 40644 56652 40646 56672
rect 40590 56616 40646 56652
rect 40682 56228 40738 56264
rect 40682 56208 40684 56228
rect 40684 56208 40736 56228
rect 40736 56208 40738 56228
rect 41050 56208 41106 56264
rect 41142 55800 41198 55856
rect 41694 55800 41750 55856
rect 41878 56344 41934 56400
rect 42338 56480 42394 56536
rect 42798 55936 42854 55992
rect 43350 55820 43406 55856
rect 43350 55800 43352 55820
rect 43352 55800 43404 55820
rect 43404 55800 43406 55820
rect 45650 56888 45706 56944
rect 45466 56652 45468 56672
rect 45468 56652 45520 56672
rect 45520 56652 45522 56672
rect 45466 56616 45522 56652
rect 45558 56244 45560 56264
rect 45560 56244 45612 56264
rect 45612 56244 45614 56264
rect 45558 56208 45614 56244
rect 44546 55392 44602 55448
rect 44730 55412 44786 55448
rect 46938 56480 46994 56536
rect 46110 56344 46166 56400
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 44730 55392 44732 55412
rect 44732 55392 44784 55412
rect 44784 55392 44786 55412
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
<< metal3 >>
rect 27521 57762 27587 57765
rect 28165 57762 28231 57765
rect 27521 57760 28231 57762
rect 27521 57704 27526 57760
rect 27582 57704 28170 57760
rect 28226 57704 28231 57760
rect 27521 57702 28231 57704
rect 27521 57699 27587 57702
rect 28165 57699 28231 57702
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 6361 57490 6427 57493
rect 27981 57490 28047 57493
rect 6361 57488 28047 57490
rect 6361 57432 6366 57488
rect 6422 57432 27986 57488
rect 28042 57432 28047 57488
rect 6361 57430 28047 57432
rect 6361 57427 6427 57430
rect 27981 57427 28047 57430
rect 11881 57354 11947 57357
rect 27705 57354 27771 57357
rect 11881 57352 27771 57354
rect 11881 57296 11886 57352
rect 11942 57296 27710 57352
rect 27766 57296 27771 57352
rect 11881 57294 27771 57296
rect 11881 57291 11947 57294
rect 27705 57291 27771 57294
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 20713 56946 20779 56949
rect 27429 56946 27495 56949
rect 20713 56944 27495 56946
rect 20713 56888 20718 56944
rect 20774 56888 27434 56944
rect 27490 56888 27495 56944
rect 20713 56886 27495 56888
rect 20713 56883 20779 56886
rect 27429 56883 27495 56886
rect 40033 56946 40099 56949
rect 45645 56946 45711 56949
rect 40033 56944 45711 56946
rect 40033 56888 40038 56944
rect 40094 56888 45650 56944
rect 45706 56888 45711 56944
rect 40033 56886 45711 56888
rect 40033 56883 40099 56886
rect 45645 56883 45711 56886
rect 27521 56810 27587 56813
rect 30005 56810 30071 56813
rect 27521 56808 30071 56810
rect 27521 56752 27526 56808
rect 27582 56752 30010 56808
rect 30066 56752 30071 56808
rect 27521 56750 30071 56752
rect 27521 56747 27587 56750
rect 30005 56747 30071 56750
rect 27705 56674 27771 56677
rect 29821 56674 29887 56677
rect 27705 56672 29887 56674
rect 27705 56616 27710 56672
rect 27766 56616 29826 56672
rect 29882 56616 29887 56672
rect 27705 56614 29887 56616
rect 27705 56611 27771 56614
rect 29821 56611 29887 56614
rect 40585 56674 40651 56677
rect 45461 56674 45527 56677
rect 40585 56672 45527 56674
rect 40585 56616 40590 56672
rect 40646 56616 45466 56672
rect 45522 56616 45527 56672
rect 40585 56614 45527 56616
rect 40585 56611 40651 56614
rect 45461 56611 45527 56614
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 29821 56538 29887 56541
rect 36077 56538 36143 56541
rect 29821 56536 36143 56538
rect 29821 56480 29826 56536
rect 29882 56480 36082 56536
rect 36138 56480 36143 56536
rect 29821 56478 36143 56480
rect 29821 56475 29887 56478
rect 36077 56475 36143 56478
rect 42333 56538 42399 56541
rect 46933 56538 46999 56541
rect 42333 56536 46999 56538
rect 42333 56480 42338 56536
rect 42394 56480 46938 56536
rect 46994 56480 46999 56536
rect 42333 56478 46999 56480
rect 42333 56475 42399 56478
rect 46933 56475 46999 56478
rect 29361 56402 29427 56405
rect 37365 56402 37431 56405
rect 29361 56400 37431 56402
rect 29361 56344 29366 56400
rect 29422 56344 37370 56400
rect 37426 56344 37431 56400
rect 29361 56342 37431 56344
rect 29361 56339 29427 56342
rect 37365 56339 37431 56342
rect 41873 56402 41939 56405
rect 46105 56402 46171 56405
rect 41873 56400 46171 56402
rect 41873 56344 41878 56400
rect 41934 56344 46110 56400
rect 46166 56344 46171 56400
rect 41873 56342 46171 56344
rect 41873 56339 41939 56342
rect 46105 56339 46171 56342
rect 26877 56266 26943 56269
rect 40677 56266 40743 56269
rect 26877 56264 40743 56266
rect 26877 56208 26882 56264
rect 26938 56208 40682 56264
rect 40738 56208 40743 56264
rect 26877 56206 40743 56208
rect 26877 56203 26943 56206
rect 40677 56203 40743 56206
rect 41045 56266 41111 56269
rect 45553 56266 45619 56269
rect 41045 56264 45619 56266
rect 41045 56208 41050 56264
rect 41106 56208 45558 56264
rect 45614 56208 45619 56264
rect 41045 56206 45619 56208
rect 41045 56203 41111 56206
rect 45553 56203 45619 56206
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 36997 55994 37063 55997
rect 37825 55994 37891 55997
rect 42793 55994 42859 55997
rect 36997 55992 42859 55994
rect 36997 55936 37002 55992
rect 37058 55936 37830 55992
rect 37886 55936 42798 55992
rect 42854 55936 42859 55992
rect 36997 55934 42859 55936
rect 36997 55931 37063 55934
rect 37825 55931 37891 55934
rect 42793 55931 42859 55934
rect 25497 55858 25563 55861
rect 41137 55858 41203 55861
rect 25497 55856 41203 55858
rect 25497 55800 25502 55856
rect 25558 55800 41142 55856
rect 41198 55800 41203 55856
rect 25497 55798 41203 55800
rect 25497 55795 25563 55798
rect 41137 55795 41203 55798
rect 41689 55858 41755 55861
rect 43345 55858 43411 55861
rect 41689 55856 43411 55858
rect 41689 55800 41694 55856
rect 41750 55800 43350 55856
rect 43406 55800 43411 55856
rect 41689 55798 43411 55800
rect 41689 55795 41755 55798
rect 43345 55795 43411 55798
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 29821 55450 29887 55453
rect 32949 55450 33015 55453
rect 29821 55448 33015 55450
rect 29821 55392 29826 55448
rect 29882 55392 32954 55448
rect 33010 55392 33015 55448
rect 29821 55390 33015 55392
rect 29821 55387 29887 55390
rect 32949 55387 33015 55390
rect 38009 55450 38075 55453
rect 44541 55450 44607 55453
rect 44725 55450 44791 55453
rect 38009 55448 44791 55450
rect 38009 55392 38014 55448
rect 38070 55392 44546 55448
rect 44602 55392 44730 55448
rect 44786 55392 44791 55448
rect 38009 55390 44791 55392
rect 38009 55387 38075 55390
rect 44541 55387 44607 55390
rect 44725 55387 44791 55390
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26312 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1666464484
transform -1 0 26404 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1666464484
transform 1 0 30636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1666464484
transform 1 0 31556 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1666464484
transform 1 0 25024 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1666464484
transform 1 0 24932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A_N
timestamp 1666464484
transform 1 0 36984 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B
timestamp 1666464484
transform 1 0 36432 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__B1
timestamp 1666464484
transform -1 0 29440 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A_N
timestamp 1666464484
transform 1 0 46276 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__B1
timestamp 1666464484
transform 1 0 39284 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B1
timestamp 1666464484
transform -1 0 28152 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1666464484
transform 1 0 35880 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__B2
timestamp 1666464484
transform 1 0 32476 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A2
timestamp 1666464484
transform -1 0 28520 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1666464484
transform 1 0 42780 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A2
timestamp 1666464484
transform -1 0 40848 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1666464484
transform 1 0 23000 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1666464484
transform -1 0 20884 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A2
timestamp 1666464484
transform -1 0 35236 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A2
timestamp 1666464484
transform 1 0 39652 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A1
timestamp 1666464484
transform -1 0 33396 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A1
timestamp 1666464484
transform 1 0 41952 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1666464484
transform 1 0 25024 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1666464484
transform 1 0 23552 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A1
timestamp 1666464484
transform 1 0 32476 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1666464484
transform 1 0 34500 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B1
timestamp 1666464484
transform -1 0 30636 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A1
timestamp 1666464484
transform -1 0 31280 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__B1
timestamp 1666464484
transform 1 0 40388 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A1
timestamp 1666464484
transform 1 0 41400 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A
timestamp 1666464484
transform 1 0 22080 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1666464484
transform 1 0 23460 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1666464484
transform 1 0 31096 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A2
timestamp 1666464484
transform 1 0 36064 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A2
timestamp 1666464484
transform 1 0 36616 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A1
timestamp 1666464484
transform -1 0 30084 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__C1
timestamp 1666464484
transform 1 0 27692 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 3680 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 28704 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 29900 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 32108 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 34132 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 35236 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 37720 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 38824 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666464484
transform -1 0 40020 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666464484
transform -1 0 46276 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666464484
transform -1 0 45724 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1666464484
transform -1 0 43884 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1666464484
transform -1 0 44712 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1666464484
transform -1 0 47104 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1666464484
transform -1 0 48024 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1666464484
transform -1 0 49404 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1666464484
transform -1 0 51244 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1666464484
transform -1 0 51796 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1666464484
transform -1 0 52532 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1666464484
transform -1 0 54004 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1666464484
transform -1 0 55292 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output22_A
timestamp 1666464484
transform 1 0 6256 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1666464484
transform 1 0 11040 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16
timestamp 1666464484
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31
timestamp 1666464484
transform 1 0 3956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1666464484
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46
timestamp 1666464484
transform 1 0 5336 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1666464484
transform 1 0 6440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61
timestamp 1666464484
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73
timestamp 1666464484
transform 1 0 7820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 1666464484
transform 1 0 8096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_88
timestamp 1666464484
transform 1 0 9200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1666464484
transform 1 0 9476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1666464484
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1666464484
transform 1 0 10580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_106
timestamp 1666464484
transform 1 0 10856 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_111
timestamp 1666464484
transform 1 0 11316 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_118
timestamp 1666464484
transform 1 0 11960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_121
timestamp 1666464484
transform 1 0 12236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_126
timestamp 1666464484
transform 1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_133
timestamp 1666464484
transform 1 0 13340 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_136
timestamp 1666464484
transform 1 0 13616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_148
timestamp 1666464484
transform 1 0 14720 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1666464484
transform 1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1666464484
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_163
timestamp 1666464484
transform 1 0 16100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1666464484
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_171
timestamp 1666464484
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1666464484
transform 1 0 17480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_186
timestamp 1666464484
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_201
timestamp 1666464484
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_208
timestamp 1666464484
transform 1 0 20240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_211
timestamp 1666464484
transform 1 0 20516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_216
timestamp 1666464484
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_223
timestamp 1666464484
transform 1 0 21620 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_226
timestamp 1666464484
transform 1 0 21896 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_231
timestamp 1666464484
transform 1 0 22356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_238
timestamp 1666464484
transform 1 0 23000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_241
timestamp 1666464484
transform 1 0 23276 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_246
timestamp 1666464484
transform 1 0 23736 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_256
timestamp 1666464484
transform 1 0 24656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_261
timestamp 1666464484
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_268
timestamp 1666464484
transform 1 0 25760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1666464484
transform 1 0 26036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1666464484
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_283
timestamp 1666464484
transform 1 0 27140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_286
timestamp 1666464484
transform 1 0 27416 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1666464484
transform 1 0 27876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_298
timestamp 1666464484
transform 1 0 28520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_301
timestamp 1666464484
transform 1 0 28796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_306
timestamp 1666464484
transform 1 0 29256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_313
timestamp 1666464484
transform 1 0 29900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_316
timestamp 1666464484
transform 1 0 30176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_320 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_324 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30912 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_331
timestamp 1666464484
transform 1 0 31556 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_336
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_343
timestamp 1666464484
transform 1 0 32660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_346
timestamp 1666464484
transform 1 0 32936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_351
timestamp 1666464484
transform 1 0 33396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_358
timestamp 1666464484
transform 1 0 34040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_361
timestamp 1666464484
transform 1 0 34316 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_366
timestamp 1666464484
transform 1 0 34776 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_373
timestamp 1666464484
transform 1 0 35420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_376
timestamp 1666464484
transform 1 0 35696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_381
timestamp 1666464484
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_388
timestamp 1666464484
transform 1 0 36800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_391
timestamp 1666464484
transform 1 0 37076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1666464484
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_403
timestamp 1666464484
transform 1 0 38180 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_406
timestamp 1666464484
transform 1 0 38456 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_411
timestamp 1666464484
transform 1 0 38916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1666464484
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1666464484
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_426
timestamp 1666464484
transform 1 0 40296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_433
timestamp 1666464484
transform 1 0 40940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_436
timestamp 1666464484
transform 1 0 41216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_441
timestamp 1666464484
transform 1 0 41676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_448
timestamp 1666464484
transform 1 0 42320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_451
timestamp 1666464484
transform 1 0 42596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_456
timestamp 1666464484
transform 1 0 43056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_463
timestamp 1666464484
transform 1 0 43700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_466
timestamp 1666464484
transform 1 0 43976 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1666464484
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_478
timestamp 1666464484
transform 1 0 45080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_481
timestamp 1666464484
transform 1 0 45356 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1666464484
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_493
timestamp 1666464484
transform 1 0 46460 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_496
timestamp 1666464484
transform 1 0 46736 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_501
timestamp 1666464484
transform 1 0 47196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_508
timestamp 1666464484
transform 1 0 47840 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_511
timestamp 1666464484
transform 1 0 48116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_516
timestamp 1666464484
transform 1 0 48576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_523
timestamp 1666464484
transform 1 0 49220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_526
timestamp 1666464484
transform 1 0 49496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_531
timestamp 1666464484
transform 1 0 49956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_538
timestamp 1666464484
transform 1 0 50600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_541
timestamp 1666464484
transform 1 0 50876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_546
timestamp 1666464484
transform 1 0 51336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_553
timestamp 1666464484
transform 1 0 51980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_556
timestamp 1666464484
transform 1 0 52256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_561
timestamp 1666464484
transform 1 0 52716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_568
timestamp 1666464484
transform 1 0 53360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_571
timestamp 1666464484
transform 1 0 53636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_576 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 54096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_584
timestamp 1666464484
transform 1 0 54832 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_586
timestamp 1666464484
transform 1 0 55016 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_598
timestamp 1666464484
transform 1 0 56120 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1666464484
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_613
timestamp 1666464484
transform 1 0 57500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_616
timestamp 1666464484
transform 1 0 57776 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_624
timestamp 1666464484
transform 1 0 58512 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1666464484
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_43
timestamp 1666464484
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_59
timestamp 1666464484
transform 1 0 6532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_61
timestamp 1666464484
transform 1 0 6716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1666464484
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_77
timestamp 1666464484
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_88
timestamp 1666464484
transform 1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_91
timestamp 1666464484
transform 1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_97
timestamp 1666464484
transform 1 0 10028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_104
timestamp 1666464484
transform 1 0 10672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1666464484
transform 1 0 11960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_121
timestamp 1666464484
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_127
timestamp 1666464484
transform 1 0 12788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_134
timestamp 1666464484
transform 1 0 13432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1666464484
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_148
timestamp 1666464484
transform 1 0 14720 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_151
timestamp 1666464484
transform 1 0 14996 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_157
timestamp 1666464484
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1666464484
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_171
timestamp 1666464484
transform 1 0 16836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_178
timestamp 1666464484
transform 1 0 17480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1666464484
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_194
timestamp 1666464484
transform 1 0 18952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1666464484
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_208
timestamp 1666464484
transform 1 0 20240 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_211
timestamp 1666464484
transform 1 0 20516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_217
timestamp 1666464484
transform 1 0 21068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_224
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_231
timestamp 1666464484
transform 1 0 22356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_238
timestamp 1666464484
transform 1 0 23000 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_241
timestamp 1666464484
transform 1 0 23276 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_268
timestamp 1666464484
transform 1 0 25760 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_271
timestamp 1666464484
transform 1 0 26036 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_298
timestamp 1666464484
transform 1 0 28520 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_301
timestamp 1666464484
transform 1 0 28796 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_328
timestamp 1666464484
transform 1 0 31280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_331
timestamp 1666464484
transform 1 0 31556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_354
timestamp 1666464484
transform 1 0 33672 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_361
timestamp 1666464484
transform 1 0 34316 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_384
timestamp 1666464484
transform 1 0 36432 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_391
timestamp 1666464484
transform 1 0 37076 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_414
timestamp 1666464484
transform 1 0 39192 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_421
timestamp 1666464484
transform 1 0 39836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_426
timestamp 1666464484
transform 1 0 40296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_433
timestamp 1666464484
transform 1 0 40940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_440
timestamp 1666464484
transform 1 0 41584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_447
timestamp 1666464484
transform 1 0 42228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_451
timestamp 1666464484
transform 1 0 42596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_456
timestamp 1666464484
transform 1 0 43056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_463
timestamp 1666464484
transform 1 0 43700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_470
timestamp 1666464484
transform 1 0 44344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_477
timestamp 1666464484
transform 1 0 44988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_481
timestamp 1666464484
transform 1 0 45356 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_486
timestamp 1666464484
transform 1 0 45816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_493
timestamp 1666464484
transform 1 0 46460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1666464484
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_507
timestamp 1666464484
transform 1 0 47748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_511
timestamp 1666464484
transform 1 0 48116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_516
timestamp 1666464484
transform 1 0 48576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_523
timestamp 1666464484
transform 1 0 49220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_530
timestamp 1666464484
transform 1 0 49864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_537
timestamp 1666464484
transform 1 0 50508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_541
timestamp 1666464484
transform 1 0 50876 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_546
timestamp 1666464484
transform 1 0 51336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_553
timestamp 1666464484
transform 1 0 51980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_560
timestamp 1666464484
transform 1 0 52624 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_567
timestamp 1666464484
transform 1 0 53268 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_571
timestamp 1666464484
transform 1 0 53636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_583
timestamp 1666464484
transform 1 0 54740 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_595
timestamp 1666464484
transform 1 0 55844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_599
timestamp 1666464484
transform 1 0 56212 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_601
timestamp 1666464484
transform 1 0 56396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_613
timestamp 1666464484
transform 1 0 57500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_16
timestamp 1666464484
transform 1 0 2576 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_28
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_40
timestamp 1666464484
transform 1 0 4784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_44
timestamp 1666464484
transform 1 0 5152 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_46
timestamp 1666464484
transform 1 0 5336 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_58
timestamp 1666464484
transform 1 0 6440 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1666464484
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_74
timestamp 1666464484
transform 1 0 7912 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_76
timestamp 1666464484
transform 1 0 8096 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_88
timestamp 1666464484
transform 1 0 9200 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_103
timestamp 1666464484
transform 1 0 10580 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_106
timestamp 1666464484
transform 1 0 10856 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_118
timestamp 1666464484
transform 1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_124
timestamp 1666464484
transform 1 0 12512 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_136
timestamp 1666464484
transform 1 0 13616 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_145
timestamp 1666464484
transform 1 0 14444 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_154
timestamp 1666464484
transform 1 0 15272 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1666464484
transform 1 0 16100 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_166
timestamp 1666464484
transform 1 0 16376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1666464484
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1666464484
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_186
timestamp 1666464484
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_193
timestamp 1666464484
transform 1 0 18860 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_196
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1666464484
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_216
timestamp 1666464484
transform 1 0 20976 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_223
timestamp 1666464484
transform 1 0 21620 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_226
timestamp 1666464484
transform 1 0 21896 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_256
timestamp 1666464484
transform 1 0 24656 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_283
timestamp 1666464484
transform 1 0 27140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_286
timestamp 1666464484
transform 1 0 27416 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_313
timestamp 1666464484
transform 1 0 29900 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_316
timestamp 1666464484
transform 1 0 30176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_341
timestamp 1666464484
transform 1 0 32476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_346
timestamp 1666464484
transform 1 0 32936 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_369
timestamp 1666464484
transform 1 0 35052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_376
timestamp 1666464484
transform 1 0 35696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_399
timestamp 1666464484
transform 1 0 37812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_406
timestamp 1666464484
transform 1 0 38456 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_411
timestamp 1666464484
transform 1 0 38916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_418
timestamp 1666464484
transform 1 0 39560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_425
timestamp 1666464484
transform 1 0 40204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_432
timestamp 1666464484
transform 1 0 40848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_436
timestamp 1666464484
transform 1 0 41216 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_441
timestamp 1666464484
transform 1 0 41676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_448
timestamp 1666464484
transform 1 0 42320 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_455
timestamp 1666464484
transform 1 0 42964 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_462
timestamp 1666464484
transform 1 0 43608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_466
timestamp 1666464484
transform 1 0 43976 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_471
timestamp 1666464484
transform 1 0 44436 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_480
timestamp 1666464484
transform 1 0 45264 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_492
timestamp 1666464484
transform 1 0 46368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_496
timestamp 1666464484
transform 1 0 46736 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_501
timestamp 1666464484
transform 1 0 47196 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_510
timestamp 1666464484
transform 1 0 48024 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_522
timestamp 1666464484
transform 1 0 49128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_526
timestamp 1666464484
transform 1 0 49496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_531
timestamp 1666464484
transform 1 0 49956 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_540
timestamp 1666464484
transform 1 0 50784 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_552
timestamp 1666464484
transform 1 0 51888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_556
timestamp 1666464484
transform 1 0 52256 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_561
timestamp 1666464484
transform 1 0 52716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_573
timestamp 1666464484
transform 1 0 53820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_586
timestamp 1666464484
transform 1 0 55016 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_598
timestamp 1666464484
transform 1 0 56120 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_610
timestamp 1666464484
transform 1 0 57224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_614
timestamp 1666464484
transform 1 0 57592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_616
timestamp 1666464484
transform 1 0 57776 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_624
timestamp 1666464484
transform 1 0 58512 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_31
timestamp 1666464484
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_43
timestamp 1666464484
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_59
timestamp 1666464484
transform 1 0 6532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_61
timestamp 1666464484
transform 1 0 6716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_73
timestamp 1666464484
transform 1 0 7820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1666464484
transform 1 0 8924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_89
timestamp 1666464484
transform 1 0 9292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_91
timestamp 1666464484
transform 1 0 9476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_103
timestamp 1666464484
transform 1 0 10580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1666464484
transform 1 0 11684 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_119
timestamp 1666464484
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_121
timestamp 1666464484
transform 1 0 12236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_133
timestamp 1666464484
transform 1 0 13340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1666464484
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_151
timestamp 1666464484
transform 1 0 14996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_163
timestamp 1666464484
transform 1 0 16100 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_178
timestamp 1666464484
transform 1 0 17480 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_192
timestamp 1666464484
transform 1 0 18768 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_201
timestamp 1666464484
transform 1 0 19596 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_208
timestamp 1666464484
transform 1 0 20240 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_211
timestamp 1666464484
transform 1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_217
timestamp 1666464484
transform 1 0 21068 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_224
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_231
timestamp 1666464484
transform 1 0 22356 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_238
timestamp 1666464484
transform 1 0 23000 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_241
timestamp 1666464484
transform 1 0 23276 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_268
timestamp 1666464484
transform 1 0 25760 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_271
timestamp 1666464484
transform 1 0 26036 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_298
timestamp 1666464484
transform 1 0 28520 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_301
timestamp 1666464484
transform 1 0 28796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_326
timestamp 1666464484
transform 1 0 31096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_331
timestamp 1666464484
transform 1 0 31556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_358
timestamp 1666464484
transform 1 0 34040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_361
timestamp 1666464484
transform 1 0 34316 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_384
timestamp 1666464484
transform 1 0 36432 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_391
timestamp 1666464484
transform 1 0 37076 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_396
timestamp 1666464484
transform 1 0 37536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1666464484
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_410
timestamp 1666464484
transform 1 0 38824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_417
timestamp 1666464484
transform 1 0 39468 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_421
timestamp 1666464484
transform 1 0 39836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_426
timestamp 1666464484
transform 1 0 40296 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_433
timestamp 1666464484
transform 1 0 40940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_445
timestamp 1666464484
transform 1 0 42044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_449
timestamp 1666464484
transform 1 0 42412 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_451
timestamp 1666464484
transform 1 0 42596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_463
timestamp 1666464484
transform 1 0 43700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_475
timestamp 1666464484
transform 1 0 44804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_479
timestamp 1666464484
transform 1 0 45172 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_481
timestamp 1666464484
transform 1 0 45356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_493
timestamp 1666464484
transform 1 0 46460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_505
timestamp 1666464484
transform 1 0 47564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_509
timestamp 1666464484
transform 1 0 47932 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_511
timestamp 1666464484
transform 1 0 48116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_523
timestamp 1666464484
transform 1 0 49220 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_535
timestamp 1666464484
transform 1 0 50324 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_539
timestamp 1666464484
transform 1 0 50692 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1666464484
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_553
timestamp 1666464484
transform 1 0 51980 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_565
timestamp 1666464484
transform 1 0 53084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_569
timestamp 1666464484
transform 1 0 53452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_571
timestamp 1666464484
transform 1 0 53636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_583
timestamp 1666464484
transform 1 0 54740 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_595
timestamp 1666464484
transform 1 0 55844 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_599
timestamp 1666464484
transform 1 0 56212 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_601
timestamp 1666464484
transform 1 0 56396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_613
timestamp 1666464484
transform 1 0 57500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_16
timestamp 1666464484
transform 1 0 2576 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_28
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_40
timestamp 1666464484
transform 1 0 4784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_44
timestamp 1666464484
transform 1 0 5152 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_46
timestamp 1666464484
transform 1 0 5336 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_58
timestamp 1666464484
transform 1 0 6440 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_70
timestamp 1666464484
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_74
timestamp 1666464484
transform 1 0 7912 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_76
timestamp 1666464484
transform 1 0 8096 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_88
timestamp 1666464484
transform 1 0 9200 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_100
timestamp 1666464484
transform 1 0 10304 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_104
timestamp 1666464484
transform 1 0 10672 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_106
timestamp 1666464484
transform 1 0 10856 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_118
timestamp 1666464484
transform 1 0 11960 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_130
timestamp 1666464484
transform 1 0 13064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_134
timestamp 1666464484
transform 1 0 13432 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_136
timestamp 1666464484
transform 1 0 13616 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_148
timestamp 1666464484
transform 1 0 14720 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_160
timestamp 1666464484
transform 1 0 15824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_164
timestamp 1666464484
transform 1 0 16192 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_166
timestamp 1666464484
transform 1 0 16376 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_178
timestamp 1666464484
transform 1 0 17480 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_190
timestamp 1666464484
transform 1 0 18584 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_194
timestamp 1666464484
transform 1 0 18952 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_196
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_208
timestamp 1666464484
transform 1 0 20240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_212
timestamp 1666464484
transform 1 0 20608 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_216
timestamp 1666464484
transform 1 0 20976 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_223
timestamp 1666464484
transform 1 0 21620 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_226
timestamp 1666464484
transform 1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_232
timestamp 1666464484
transform 1 0 22448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_239
timestamp 1666464484
transform 1 0 23092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_246
timestamp 1666464484
transform 1 0 23736 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_256
timestamp 1666464484
transform 1 0 24656 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_283
timestamp 1666464484
transform 1 0 27140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_286
timestamp 1666464484
transform 1 0 27416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_316
timestamp 1666464484
transform 1 0 30176 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_339
timestamp 1666464484
transform 1 0 32292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_346
timestamp 1666464484
transform 1 0 32936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_369
timestamp 1666464484
transform 1 0 35052 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_376
timestamp 1666464484
transform 1 0 35696 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_381
timestamp 1666464484
transform 1 0 36156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_388
timestamp 1666464484
transform 1 0 36800 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_395
timestamp 1666464484
transform 1 0 37444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_402
timestamp 1666464484
transform 1 0 38088 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_406
timestamp 1666464484
transform 1 0 38456 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_418
timestamp 1666464484
transform 1 0 39560 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_430
timestamp 1666464484
transform 1 0 40664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_434
timestamp 1666464484
transform 1 0 41032 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_436
timestamp 1666464484
transform 1 0 41216 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_448
timestamp 1666464484
transform 1 0 42320 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_460
timestamp 1666464484
transform 1 0 43424 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_464
timestamp 1666464484
transform 1 0 43792 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_466
timestamp 1666464484
transform 1 0 43976 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_478
timestamp 1666464484
transform 1 0 45080 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_490
timestamp 1666464484
transform 1 0 46184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_494
timestamp 1666464484
transform 1 0 46552 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_496
timestamp 1666464484
transform 1 0 46736 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_508
timestamp 1666464484
transform 1 0 47840 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_520
timestamp 1666464484
transform 1 0 48944 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_524
timestamp 1666464484
transform 1 0 49312 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_526
timestamp 1666464484
transform 1 0 49496 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_538
timestamp 1666464484
transform 1 0 50600 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_550
timestamp 1666464484
transform 1 0 51704 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_554
timestamp 1666464484
transform 1 0 52072 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_556
timestamp 1666464484
transform 1 0 52256 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_568
timestamp 1666464484
transform 1 0 53360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_580
timestamp 1666464484
transform 1 0 54464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_584
timestamp 1666464484
transform 1 0 54832 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_586
timestamp 1666464484
transform 1 0 55016 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_598
timestamp 1666464484
transform 1 0 56120 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_610
timestamp 1666464484
transform 1 0 57224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_614
timestamp 1666464484
transform 1 0 57592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_616
timestamp 1666464484
transform 1 0 57776 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_624
timestamp 1666464484
transform 1 0 58512 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_31
timestamp 1666464484
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_43
timestamp 1666464484
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_59
timestamp 1666464484
transform 1 0 6532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_61
timestamp 1666464484
transform 1 0 6716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_73
timestamp 1666464484
transform 1 0 7820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_85
timestamp 1666464484
transform 1 0 8924 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_89
timestamp 1666464484
transform 1 0 9292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_91
timestamp 1666464484
transform 1 0 9476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_103
timestamp 1666464484
transform 1 0 10580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_115
timestamp 1666464484
transform 1 0 11684 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_119
timestamp 1666464484
transform 1 0 12052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_121
timestamp 1666464484
transform 1 0 12236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_133
timestamp 1666464484
transform 1 0 13340 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1666464484
transform 1 0 14444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_151
timestamp 1666464484
transform 1 0 14996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_163
timestamp 1666464484
transform 1 0 16100 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_175
timestamp 1666464484
transform 1 0 17204 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_179
timestamp 1666464484
transform 1 0 17572 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_209
timestamp 1666464484
transform 1 0 20332 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_211
timestamp 1666464484
transform 1 0 20516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_231
timestamp 1666464484
transform 1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_241
timestamp 1666464484
transform 1 0 23276 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1666464484
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_251
timestamp 1666464484
transform 1 0 24196 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_258
timestamp 1666464484
transform 1 0 24840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_268
timestamp 1666464484
transform 1 0 25760 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_271
timestamp 1666464484
transform 1 0 26036 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_298
timestamp 1666464484
transform 1 0 28520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_301
timestamp 1666464484
transform 1 0 28796 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_328
timestamp 1666464484
transform 1 0 31280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_331
timestamp 1666464484
transform 1 0 31556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_354
timestamp 1666464484
transform 1 0 33672 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_361
timestamp 1666464484
transform 1 0 34316 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_384
timestamp 1666464484
transform 1 0 36432 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_391
timestamp 1666464484
transform 1 0 37076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_403
timestamp 1666464484
transform 1 0 38180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_415
timestamp 1666464484
transform 1 0 39284 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_419
timestamp 1666464484
transform 1 0 39652 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_421
timestamp 1666464484
transform 1 0 39836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_433
timestamp 1666464484
transform 1 0 40940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_445
timestamp 1666464484
transform 1 0 42044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_449
timestamp 1666464484
transform 1 0 42412 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_451
timestamp 1666464484
transform 1 0 42596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_463
timestamp 1666464484
transform 1 0 43700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_475
timestamp 1666464484
transform 1 0 44804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_479
timestamp 1666464484
transform 1 0 45172 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_481
timestamp 1666464484
transform 1 0 45356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_493
timestamp 1666464484
transform 1 0 46460 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_505
timestamp 1666464484
transform 1 0 47564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_509
timestamp 1666464484
transform 1 0 47932 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_511
timestamp 1666464484
transform 1 0 48116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_523
timestamp 1666464484
transform 1 0 49220 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_535
timestamp 1666464484
transform 1 0 50324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_539
timestamp 1666464484
transform 1 0 50692 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1666464484
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_553
timestamp 1666464484
transform 1 0 51980 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_565
timestamp 1666464484
transform 1 0 53084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_569
timestamp 1666464484
transform 1 0 53452 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_571
timestamp 1666464484
transform 1 0 53636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_583
timestamp 1666464484
transform 1 0 54740 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_595
timestamp 1666464484
transform 1 0 55844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_599
timestamp 1666464484
transform 1 0 56212 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_601
timestamp 1666464484
transform 1 0 56396 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_613
timestamp 1666464484
transform 1 0 57500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_16
timestamp 1666464484
transform 1 0 2576 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_28
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_40
timestamp 1666464484
transform 1 0 4784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_44
timestamp 1666464484
transform 1 0 5152 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_46
timestamp 1666464484
transform 1 0 5336 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_58
timestamp 1666464484
transform 1 0 6440 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_70
timestamp 1666464484
transform 1 0 7544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_74
timestamp 1666464484
transform 1 0 7912 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_76
timestamp 1666464484
transform 1 0 8096 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_88
timestamp 1666464484
transform 1 0 9200 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_100
timestamp 1666464484
transform 1 0 10304 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_104
timestamp 1666464484
transform 1 0 10672 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_106
timestamp 1666464484
transform 1 0 10856 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_118
timestamp 1666464484
transform 1 0 11960 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_130
timestamp 1666464484
transform 1 0 13064 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_134
timestamp 1666464484
transform 1 0 13432 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_136
timestamp 1666464484
transform 1 0 13616 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_148
timestamp 1666464484
transform 1 0 14720 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_160
timestamp 1666464484
transform 1 0 15824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_164
timestamp 1666464484
transform 1 0 16192 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_166
timestamp 1666464484
transform 1 0 16376 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_178
timestamp 1666464484
transform 1 0 17480 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_190
timestamp 1666464484
transform 1 0 18584 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_194
timestamp 1666464484
transform 1 0 18952 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_196
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_208
timestamp 1666464484
transform 1 0 20240 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_220
timestamp 1666464484
transform 1 0 21344 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_224
timestamp 1666464484
transform 1 0 21712 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_226
timestamp 1666464484
transform 1 0 21896 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_238
timestamp 1666464484
transform 1 0 23000 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_242
timestamp 1666464484
transform 1 0 23368 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_246
timestamp 1666464484
transform 1 0 23736 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_256
timestamp 1666464484
transform 1 0 24656 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_283
timestamp 1666464484
transform 1 0 27140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_286
timestamp 1666464484
transform 1 0 27416 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_290
timestamp 1666464484
transform 1 0 27784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_312
timestamp 1666464484
transform 1 0 29808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_316
timestamp 1666464484
transform 1 0 30176 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_343
timestamp 1666464484
transform 1 0 32660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_346
timestamp 1666464484
transform 1 0 32936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_369
timestamp 1666464484
transform 1 0 35052 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_376
timestamp 1666464484
transform 1 0 35696 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_388
timestamp 1666464484
transform 1 0 36800 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_400
timestamp 1666464484
transform 1 0 37904 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_404
timestamp 1666464484
transform 1 0 38272 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_406
timestamp 1666464484
transform 1 0 38456 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_418
timestamp 1666464484
transform 1 0 39560 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_430
timestamp 1666464484
transform 1 0 40664 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_434
timestamp 1666464484
transform 1 0 41032 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_436
timestamp 1666464484
transform 1 0 41216 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_448
timestamp 1666464484
transform 1 0 42320 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_460
timestamp 1666464484
transform 1 0 43424 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_464
timestamp 1666464484
transform 1 0 43792 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_466
timestamp 1666464484
transform 1 0 43976 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_478
timestamp 1666464484
transform 1 0 45080 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_490
timestamp 1666464484
transform 1 0 46184 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_494
timestamp 1666464484
transform 1 0 46552 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_496
timestamp 1666464484
transform 1 0 46736 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_508
timestamp 1666464484
transform 1 0 47840 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_520
timestamp 1666464484
transform 1 0 48944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_524
timestamp 1666464484
transform 1 0 49312 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_526
timestamp 1666464484
transform 1 0 49496 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_538
timestamp 1666464484
transform 1 0 50600 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_550
timestamp 1666464484
transform 1 0 51704 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_554
timestamp 1666464484
transform 1 0 52072 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_556
timestamp 1666464484
transform 1 0 52256 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_568
timestamp 1666464484
transform 1 0 53360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_580
timestamp 1666464484
transform 1 0 54464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_584
timestamp 1666464484
transform 1 0 54832 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_586
timestamp 1666464484
transform 1 0 55016 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_598
timestamp 1666464484
transform 1 0 56120 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_610
timestamp 1666464484
transform 1 0 57224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_614
timestamp 1666464484
transform 1 0 57592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_616
timestamp 1666464484
transform 1 0 57776 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_624
timestamp 1666464484
transform 1 0 58512 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_31
timestamp 1666464484
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_43
timestamp 1666464484
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_59
timestamp 1666464484
transform 1 0 6532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_61
timestamp 1666464484
transform 1 0 6716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_73
timestamp 1666464484
transform 1 0 7820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_85
timestamp 1666464484
transform 1 0 8924 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_89
timestamp 1666464484
transform 1 0 9292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_91
timestamp 1666464484
transform 1 0 9476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_103
timestamp 1666464484
transform 1 0 10580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_115
timestamp 1666464484
transform 1 0 11684 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_119
timestamp 1666464484
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_121
timestamp 1666464484
transform 1 0 12236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_133
timestamp 1666464484
transform 1 0 13340 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1666464484
transform 1 0 14444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_151
timestamp 1666464484
transform 1 0 14996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_163
timestamp 1666464484
transform 1 0 16100 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_175
timestamp 1666464484
transform 1 0 17204 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_179
timestamp 1666464484
transform 1 0 17572 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_209
timestamp 1666464484
transform 1 0 20332 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_211
timestamp 1666464484
transform 1 0 20516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_235
timestamp 1666464484
transform 1 0 22724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_239
timestamp 1666464484
transform 1 0 23092 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_241
timestamp 1666464484
transform 1 0 23276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_253
timestamp 1666464484
transform 1 0 24380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_268
timestamp 1666464484
transform 1 0 25760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_271
timestamp 1666464484
transform 1 0 26036 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_298
timestamp 1666464484
transform 1 0 28520 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_301
timestamp 1666464484
transform 1 0 28796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_305
timestamp 1666464484
transform 1 0 29164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_327
timestamp 1666464484
transform 1 0 31188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_331
timestamp 1666464484
transform 1 0 31556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_339
timestamp 1666464484
transform 1 0 32292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_346
timestamp 1666464484
transform 1 0 32936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_353
timestamp 1666464484
transform 1 0 33580 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_359
timestamp 1666464484
transform 1 0 34132 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_361
timestamp 1666464484
transform 1 0 34316 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_366
timestamp 1666464484
transform 1 0 34776 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_378
timestamp 1666464484
transform 1 0 35880 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_391
timestamp 1666464484
transform 1 0 37076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_403
timestamp 1666464484
transform 1 0 38180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_415
timestamp 1666464484
transform 1 0 39284 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_419
timestamp 1666464484
transform 1 0 39652 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_421
timestamp 1666464484
transform 1 0 39836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_433
timestamp 1666464484
transform 1 0 40940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_445
timestamp 1666464484
transform 1 0 42044 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_449
timestamp 1666464484
transform 1 0 42412 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_451
timestamp 1666464484
transform 1 0 42596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_463
timestamp 1666464484
transform 1 0 43700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_475
timestamp 1666464484
transform 1 0 44804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_479
timestamp 1666464484
transform 1 0 45172 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_481
timestamp 1666464484
transform 1 0 45356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_493
timestamp 1666464484
transform 1 0 46460 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1666464484
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_509
timestamp 1666464484
transform 1 0 47932 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_511
timestamp 1666464484
transform 1 0 48116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_523
timestamp 1666464484
transform 1 0 49220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_535
timestamp 1666464484
transform 1 0 50324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_539
timestamp 1666464484
transform 1 0 50692 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1666464484
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_553
timestamp 1666464484
transform 1 0 51980 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_565
timestamp 1666464484
transform 1 0 53084 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_569
timestamp 1666464484
transform 1 0 53452 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_571
timestamp 1666464484
transform 1 0 53636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_583
timestamp 1666464484
transform 1 0 54740 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_595
timestamp 1666464484
transform 1 0 55844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_599
timestamp 1666464484
transform 1 0 56212 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_601
timestamp 1666464484
transform 1 0 56396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_613
timestamp 1666464484
transform 1 0 57500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_16
timestamp 1666464484
transform 1 0 2576 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_28
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_40
timestamp 1666464484
transform 1 0 4784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_44
timestamp 1666464484
transform 1 0 5152 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_46
timestamp 1666464484
transform 1 0 5336 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_58
timestamp 1666464484
transform 1 0 6440 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_70
timestamp 1666464484
transform 1 0 7544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_74
timestamp 1666464484
transform 1 0 7912 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_76
timestamp 1666464484
transform 1 0 8096 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_88
timestamp 1666464484
transform 1 0 9200 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_100
timestamp 1666464484
transform 1 0 10304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_104
timestamp 1666464484
transform 1 0 10672 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_106
timestamp 1666464484
transform 1 0 10856 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_118
timestamp 1666464484
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_130
timestamp 1666464484
transform 1 0 13064 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_134
timestamp 1666464484
transform 1 0 13432 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_136
timestamp 1666464484
transform 1 0 13616 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_148
timestamp 1666464484
transform 1 0 14720 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_160
timestamp 1666464484
transform 1 0 15824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_164
timestamp 1666464484
transform 1 0 16192 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_166
timestamp 1666464484
transform 1 0 16376 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_178
timestamp 1666464484
transform 1 0 17480 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_190
timestamp 1666464484
transform 1 0 18584 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_194
timestamp 1666464484
transform 1 0 18952 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_196
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_208
timestamp 1666464484
transform 1 0 20240 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_220
timestamp 1666464484
transform 1 0 21344 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_224
timestamp 1666464484
transform 1 0 21712 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_226
timestamp 1666464484
transform 1 0 21896 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_238
timestamp 1666464484
transform 1 0 23000 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_250
timestamp 1666464484
transform 1 0 24104 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_254
timestamp 1666464484
transform 1 0 24472 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_256
timestamp 1666464484
transform 1 0 24656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_262
timestamp 1666464484
transform 1 0 25208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_269
timestamp 1666464484
transform 1 0 25852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_276
timestamp 1666464484
transform 1 0 26496 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_283
timestamp 1666464484
transform 1 0 27140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_286
timestamp 1666464484
transform 1 0 27416 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_291
timestamp 1666464484
transform 1 0 27876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_298
timestamp 1666464484
transform 1 0 28520 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_305
timestamp 1666464484
transform 1 0 29164 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_312
timestamp 1666464484
transform 1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_316
timestamp 1666464484
transform 1 0 30176 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_322
timestamp 1666464484
transform 1 0 30728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_329
timestamp 1666464484
transform 1 0 31372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_336
timestamp 1666464484
transform 1 0 32016 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_343
timestamp 1666464484
transform 1 0 32660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_346
timestamp 1666464484
transform 1 0 32936 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_351
timestamp 1666464484
transform 1 0 33396 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_358
timestamp 1666464484
transform 1 0 34040 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_370
timestamp 1666464484
transform 1 0 35144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_374
timestamp 1666464484
transform 1 0 35512 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_376
timestamp 1666464484
transform 1 0 35696 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_388
timestamp 1666464484
transform 1 0 36800 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_400
timestamp 1666464484
transform 1 0 37904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_404
timestamp 1666464484
transform 1 0 38272 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_406
timestamp 1666464484
transform 1 0 38456 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_418
timestamp 1666464484
transform 1 0 39560 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_430
timestamp 1666464484
transform 1 0 40664 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_434
timestamp 1666464484
transform 1 0 41032 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_436
timestamp 1666464484
transform 1 0 41216 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_448
timestamp 1666464484
transform 1 0 42320 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_460
timestamp 1666464484
transform 1 0 43424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_464
timestamp 1666464484
transform 1 0 43792 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_466
timestamp 1666464484
transform 1 0 43976 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_478
timestamp 1666464484
transform 1 0 45080 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_490
timestamp 1666464484
transform 1 0 46184 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_494
timestamp 1666464484
transform 1 0 46552 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_496
timestamp 1666464484
transform 1 0 46736 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_508
timestamp 1666464484
transform 1 0 47840 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_520
timestamp 1666464484
transform 1 0 48944 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_524
timestamp 1666464484
transform 1 0 49312 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_526
timestamp 1666464484
transform 1 0 49496 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_538
timestamp 1666464484
transform 1 0 50600 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_550
timestamp 1666464484
transform 1 0 51704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_554
timestamp 1666464484
transform 1 0 52072 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_556
timestamp 1666464484
transform 1 0 52256 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_568
timestamp 1666464484
transform 1 0 53360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_580
timestamp 1666464484
transform 1 0 54464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_584
timestamp 1666464484
transform 1 0 54832 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_586
timestamp 1666464484
transform 1 0 55016 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_598
timestamp 1666464484
transform 1 0 56120 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_610
timestamp 1666464484
transform 1 0 57224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_614
timestamp 1666464484
transform 1 0 57592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_616
timestamp 1666464484
transform 1 0 57776 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_624
timestamp 1666464484
transform 1 0 58512 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_31
timestamp 1666464484
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_43
timestamp 1666464484
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_59
timestamp 1666464484
transform 1 0 6532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_61
timestamp 1666464484
transform 1 0 6716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_73
timestamp 1666464484
transform 1 0 7820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_85
timestamp 1666464484
transform 1 0 8924 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_89
timestamp 1666464484
transform 1 0 9292 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_91
timestamp 1666464484
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_103
timestamp 1666464484
transform 1 0 10580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_115
timestamp 1666464484
transform 1 0 11684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_119
timestamp 1666464484
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_121
timestamp 1666464484
transform 1 0 12236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_133
timestamp 1666464484
transform 1 0 13340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_145
timestamp 1666464484
transform 1 0 14444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_151
timestamp 1666464484
transform 1 0 14996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_163
timestamp 1666464484
transform 1 0 16100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_175
timestamp 1666464484
transform 1 0 17204 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_179
timestamp 1666464484
transform 1 0 17572 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_205
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_209
timestamp 1666464484
transform 1 0 20332 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_211
timestamp 1666464484
transform 1 0 20516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_235
timestamp 1666464484
transform 1 0 22724 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_239
timestamp 1666464484
transform 1 0 23092 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_241
timestamp 1666464484
transform 1 0 23276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1666464484
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_265
timestamp 1666464484
transform 1 0 25484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_269
timestamp 1666464484
transform 1 0 25852 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_271
timestamp 1666464484
transform 1 0 26036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_283
timestamp 1666464484
transform 1 0 27140 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_288
timestamp 1666464484
transform 1 0 27600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1666464484
transform 1 0 28244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_299
timestamp 1666464484
transform 1 0 28612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_301
timestamp 1666464484
transform 1 0 28796 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_307
timestamp 1666464484
transform 1 0 29348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_311
timestamp 1666464484
transform 1 0 29716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_318
timestamp 1666464484
transform 1 0 30360 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_325
timestamp 1666464484
transform 1 0 31004 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_329
timestamp 1666464484
transform 1 0 31372 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1666464484
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1666464484
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_339
timestamp 1666464484
transform 1 0 32292 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_346
timestamp 1666464484
transform 1 0 32936 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_358
timestamp 1666464484
transform 1 0 34040 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1666464484
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1666464484
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_385
timestamp 1666464484
transform 1 0 36524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_389
timestamp 1666464484
transform 1 0 36892 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_391
timestamp 1666464484
transform 1 0 37076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_403
timestamp 1666464484
transform 1 0 38180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_415
timestamp 1666464484
transform 1 0 39284 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_419
timestamp 1666464484
transform 1 0 39652 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_421
timestamp 1666464484
transform 1 0 39836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_433
timestamp 1666464484
transform 1 0 40940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_445
timestamp 1666464484
transform 1 0 42044 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_449
timestamp 1666464484
transform 1 0 42412 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_451
timestamp 1666464484
transform 1 0 42596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_463
timestamp 1666464484
transform 1 0 43700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_475
timestamp 1666464484
transform 1 0 44804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_479
timestamp 1666464484
transform 1 0 45172 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_481
timestamp 1666464484
transform 1 0 45356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_493
timestamp 1666464484
transform 1 0 46460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1666464484
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_509
timestamp 1666464484
transform 1 0 47932 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_511
timestamp 1666464484
transform 1 0 48116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_523
timestamp 1666464484
transform 1 0 49220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_535
timestamp 1666464484
transform 1 0 50324 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_539
timestamp 1666464484
transform 1 0 50692 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1666464484
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_553
timestamp 1666464484
transform 1 0 51980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_565
timestamp 1666464484
transform 1 0 53084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_569
timestamp 1666464484
transform 1 0 53452 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_571
timestamp 1666464484
transform 1 0 53636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_583
timestamp 1666464484
transform 1 0 54740 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_595
timestamp 1666464484
transform 1 0 55844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_599
timestamp 1666464484
transform 1 0 56212 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_601
timestamp 1666464484
transform 1 0 56396 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_613
timestamp 1666464484
transform 1 0 57500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_16
timestamp 1666464484
transform 1 0 2576 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_28
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_40
timestamp 1666464484
transform 1 0 4784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_44
timestamp 1666464484
transform 1 0 5152 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_46
timestamp 1666464484
transform 1 0 5336 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_58
timestamp 1666464484
transform 1 0 6440 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_70
timestamp 1666464484
transform 1 0 7544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_74
timestamp 1666464484
transform 1 0 7912 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_76
timestamp 1666464484
transform 1 0 8096 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_88
timestamp 1666464484
transform 1 0 9200 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1666464484
transform 1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_104
timestamp 1666464484
transform 1 0 10672 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_106
timestamp 1666464484
transform 1 0 10856 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_118
timestamp 1666464484
transform 1 0 11960 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_130
timestamp 1666464484
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_134
timestamp 1666464484
transform 1 0 13432 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_136
timestamp 1666464484
transform 1 0 13616 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_148
timestamp 1666464484
transform 1 0 14720 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_160
timestamp 1666464484
transform 1 0 15824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_164
timestamp 1666464484
transform 1 0 16192 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_166
timestamp 1666464484
transform 1 0 16376 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_178
timestamp 1666464484
transform 1 0 17480 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_190
timestamp 1666464484
transform 1 0 18584 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_194
timestamp 1666464484
transform 1 0 18952 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_196
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_208
timestamp 1666464484
transform 1 0 20240 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_220
timestamp 1666464484
transform 1 0 21344 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_224
timestamp 1666464484
transform 1 0 21712 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_226
timestamp 1666464484
transform 1 0 21896 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_238
timestamp 1666464484
transform 1 0 23000 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_250
timestamp 1666464484
transform 1 0 24104 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_254
timestamp 1666464484
transform 1 0 24472 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_256
timestamp 1666464484
transform 1 0 24656 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_268
timestamp 1666464484
transform 1 0 25760 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_280
timestamp 1666464484
transform 1 0 26864 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_284
timestamp 1666464484
transform 1 0 27232 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_286
timestamp 1666464484
transform 1 0 27416 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_298
timestamp 1666464484
transform 1 0 28520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_306
timestamp 1666464484
transform 1 0 29256 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_310
timestamp 1666464484
transform 1 0 29624 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_314
timestamp 1666464484
transform 1 0 29992 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_316
timestamp 1666464484
transform 1 0 30176 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_320
timestamp 1666464484
transform 1 0 30544 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_323
timestamp 1666464484
transform 1 0 30820 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1666464484
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_346
timestamp 1666464484
transform 1 0 32936 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_358
timestamp 1666464484
transform 1 0 34040 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_370
timestamp 1666464484
transform 1 0 35144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_374
timestamp 1666464484
transform 1 0 35512 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_376
timestamp 1666464484
transform 1 0 35696 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_388
timestamp 1666464484
transform 1 0 36800 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_400
timestamp 1666464484
transform 1 0 37904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_404
timestamp 1666464484
transform 1 0 38272 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_406
timestamp 1666464484
transform 1 0 38456 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_418
timestamp 1666464484
transform 1 0 39560 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_430
timestamp 1666464484
transform 1 0 40664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_434
timestamp 1666464484
transform 1 0 41032 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_436
timestamp 1666464484
transform 1 0 41216 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_448
timestamp 1666464484
transform 1 0 42320 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_460
timestamp 1666464484
transform 1 0 43424 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_464
timestamp 1666464484
transform 1 0 43792 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_466
timestamp 1666464484
transform 1 0 43976 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_478
timestamp 1666464484
transform 1 0 45080 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_490
timestamp 1666464484
transform 1 0 46184 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_494
timestamp 1666464484
transform 1 0 46552 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_496
timestamp 1666464484
transform 1 0 46736 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_508
timestamp 1666464484
transform 1 0 47840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_520
timestamp 1666464484
transform 1 0 48944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_524
timestamp 1666464484
transform 1 0 49312 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_526
timestamp 1666464484
transform 1 0 49496 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_538
timestamp 1666464484
transform 1 0 50600 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_550
timestamp 1666464484
transform 1 0 51704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_554
timestamp 1666464484
transform 1 0 52072 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_556
timestamp 1666464484
transform 1 0 52256 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_568
timestamp 1666464484
transform 1 0 53360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_580
timestamp 1666464484
transform 1 0 54464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_584
timestamp 1666464484
transform 1 0 54832 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_586
timestamp 1666464484
transform 1 0 55016 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_598
timestamp 1666464484
transform 1 0 56120 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_610
timestamp 1666464484
transform 1 0 57224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_614
timestamp 1666464484
transform 1 0 57592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_616
timestamp 1666464484
transform 1 0 57776 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_624
timestamp 1666464484
transform 1 0 58512 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1666464484
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1666464484
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_59
timestamp 1666464484
transform 1 0 6532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_61
timestamp 1666464484
transform 1 0 6716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_73
timestamp 1666464484
transform 1 0 7820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1666464484
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_89
timestamp 1666464484
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_91
timestamp 1666464484
transform 1 0 9476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_103
timestamp 1666464484
transform 1 0 10580 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1666464484
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_119
timestamp 1666464484
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_121
timestamp 1666464484
transform 1 0 12236 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_133
timestamp 1666464484
transform 1 0 13340 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_145
timestamp 1666464484
transform 1 0 14444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_151
timestamp 1666464484
transform 1 0 14996 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_163
timestamp 1666464484
transform 1 0 16100 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_175
timestamp 1666464484
transform 1 0 17204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_179
timestamp 1666464484
transform 1 0 17572 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_209
timestamp 1666464484
transform 1 0 20332 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_211
timestamp 1666464484
transform 1 0 20516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_235
timestamp 1666464484
transform 1 0 22724 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_239
timestamp 1666464484
transform 1 0 23092 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_241
timestamp 1666464484
transform 1 0 23276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_253
timestamp 1666464484
transform 1 0 24380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_265
timestamp 1666464484
transform 1 0 25484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_269
timestamp 1666464484
transform 1 0 25852 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_271
timestamp 1666464484
transform 1 0 26036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_283
timestamp 1666464484
transform 1 0 27140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_295
timestamp 1666464484
transform 1 0 28244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_299
timestamp 1666464484
transform 1 0 28612 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_301
timestamp 1666464484
transform 1 0 28796 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_313
timestamp 1666464484
transform 1 0 29900 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_325
timestamp 1666464484
transform 1 0 31004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_329
timestamp 1666464484
transform 1 0 31372 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_331
timestamp 1666464484
transform 1 0 31556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_343
timestamp 1666464484
transform 1 0 32660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_355
timestamp 1666464484
transform 1 0 33764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_359
timestamp 1666464484
transform 1 0 34132 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1666464484
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1666464484
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_385
timestamp 1666464484
transform 1 0 36524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_389
timestamp 1666464484
transform 1 0 36892 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_391
timestamp 1666464484
transform 1 0 37076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_403
timestamp 1666464484
transform 1 0 38180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_415
timestamp 1666464484
transform 1 0 39284 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_419
timestamp 1666464484
transform 1 0 39652 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_421
timestamp 1666464484
transform 1 0 39836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_433
timestamp 1666464484
transform 1 0 40940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_445
timestamp 1666464484
transform 1 0 42044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_449
timestamp 1666464484
transform 1 0 42412 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_451
timestamp 1666464484
transform 1 0 42596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_463
timestamp 1666464484
transform 1 0 43700 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_475
timestamp 1666464484
transform 1 0 44804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_479
timestamp 1666464484
transform 1 0 45172 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_481
timestamp 1666464484
transform 1 0 45356 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_493
timestamp 1666464484
transform 1 0 46460 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1666464484
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_509
timestamp 1666464484
transform 1 0 47932 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_511
timestamp 1666464484
transform 1 0 48116 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_523
timestamp 1666464484
transform 1 0 49220 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_535
timestamp 1666464484
transform 1 0 50324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_539
timestamp 1666464484
transform 1 0 50692 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1666464484
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_553
timestamp 1666464484
transform 1 0 51980 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_565
timestamp 1666464484
transform 1 0 53084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_569
timestamp 1666464484
transform 1 0 53452 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_571
timestamp 1666464484
transform 1 0 53636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_583
timestamp 1666464484
transform 1 0 54740 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_595
timestamp 1666464484
transform 1 0 55844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_599
timestamp 1666464484
transform 1 0 56212 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_601
timestamp 1666464484
transform 1 0 56396 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_613
timestamp 1666464484
transform 1 0 57500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_16
timestamp 1666464484
transform 1 0 2576 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_28
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_40
timestamp 1666464484
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_44
timestamp 1666464484
transform 1 0 5152 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_46
timestamp 1666464484
transform 1 0 5336 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_58
timestamp 1666464484
transform 1 0 6440 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_70
timestamp 1666464484
transform 1 0 7544 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_74
timestamp 1666464484
transform 1 0 7912 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_76
timestamp 1666464484
transform 1 0 8096 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_88
timestamp 1666464484
transform 1 0 9200 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_100
timestamp 1666464484
transform 1 0 10304 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_104
timestamp 1666464484
transform 1 0 10672 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_106
timestamp 1666464484
transform 1 0 10856 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_118
timestamp 1666464484
transform 1 0 11960 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_130
timestamp 1666464484
transform 1 0 13064 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1666464484
transform 1 0 13432 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_136
timestamp 1666464484
transform 1 0 13616 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_148
timestamp 1666464484
transform 1 0 14720 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_160
timestamp 1666464484
transform 1 0 15824 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_164
timestamp 1666464484
transform 1 0 16192 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_166
timestamp 1666464484
transform 1 0 16376 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_178
timestamp 1666464484
transform 1 0 17480 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_190
timestamp 1666464484
transform 1 0 18584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_194
timestamp 1666464484
transform 1 0 18952 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_196
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_208
timestamp 1666464484
transform 1 0 20240 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_220
timestamp 1666464484
transform 1 0 21344 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_224
timestamp 1666464484
transform 1 0 21712 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_226
timestamp 1666464484
transform 1 0 21896 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_238
timestamp 1666464484
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_250
timestamp 1666464484
transform 1 0 24104 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_254
timestamp 1666464484
transform 1 0 24472 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_256
timestamp 1666464484
transform 1 0 24656 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_268
timestamp 1666464484
transform 1 0 25760 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_280
timestamp 1666464484
transform 1 0 26864 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_284
timestamp 1666464484
transform 1 0 27232 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_286
timestamp 1666464484
transform 1 0 27416 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_298
timestamp 1666464484
transform 1 0 28520 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_310
timestamp 1666464484
transform 1 0 29624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_314
timestamp 1666464484
transform 1 0 29992 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_316
timestamp 1666464484
transform 1 0 30176 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_328
timestamp 1666464484
transform 1 0 31280 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_340
timestamp 1666464484
transform 1 0 32384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_344
timestamp 1666464484
transform 1 0 32752 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_346
timestamp 1666464484
transform 1 0 32936 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_358
timestamp 1666464484
transform 1 0 34040 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_370
timestamp 1666464484
transform 1 0 35144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_374
timestamp 1666464484
transform 1 0 35512 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_376
timestamp 1666464484
transform 1 0 35696 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_388
timestamp 1666464484
transform 1 0 36800 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_400
timestamp 1666464484
transform 1 0 37904 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_404
timestamp 1666464484
transform 1 0 38272 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_406
timestamp 1666464484
transform 1 0 38456 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_418
timestamp 1666464484
transform 1 0 39560 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_430
timestamp 1666464484
transform 1 0 40664 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_434
timestamp 1666464484
transform 1 0 41032 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_436
timestamp 1666464484
transform 1 0 41216 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_448
timestamp 1666464484
transform 1 0 42320 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_460
timestamp 1666464484
transform 1 0 43424 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_464
timestamp 1666464484
transform 1 0 43792 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_466
timestamp 1666464484
transform 1 0 43976 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_478
timestamp 1666464484
transform 1 0 45080 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_490
timestamp 1666464484
transform 1 0 46184 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_494
timestamp 1666464484
transform 1 0 46552 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_496
timestamp 1666464484
transform 1 0 46736 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_508
timestamp 1666464484
transform 1 0 47840 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_520
timestamp 1666464484
transform 1 0 48944 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_524
timestamp 1666464484
transform 1 0 49312 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_526
timestamp 1666464484
transform 1 0 49496 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_538
timestamp 1666464484
transform 1 0 50600 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_550
timestamp 1666464484
transform 1 0 51704 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_554
timestamp 1666464484
transform 1 0 52072 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_556
timestamp 1666464484
transform 1 0 52256 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_568
timestamp 1666464484
transform 1 0 53360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_580
timestamp 1666464484
transform 1 0 54464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_584
timestamp 1666464484
transform 1 0 54832 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_586
timestamp 1666464484
transform 1 0 55016 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_598
timestamp 1666464484
transform 1 0 56120 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_610
timestamp 1666464484
transform 1 0 57224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_614
timestamp 1666464484
transform 1 0 57592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_616
timestamp 1666464484
transform 1 0 57776 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_624
timestamp 1666464484
transform 1 0 58512 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_27
timestamp 1666464484
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_31
timestamp 1666464484
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_43
timestamp 1666464484
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_55
timestamp 1666464484
transform 1 0 6164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_59
timestamp 1666464484
transform 1 0 6532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_61
timestamp 1666464484
transform 1 0 6716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_73
timestamp 1666464484
transform 1 0 7820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_85
timestamp 1666464484
transform 1 0 8924 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_89
timestamp 1666464484
transform 1 0 9292 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_91
timestamp 1666464484
transform 1 0 9476 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_103
timestamp 1666464484
transform 1 0 10580 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1666464484
transform 1 0 11684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1666464484
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_121
timestamp 1666464484
transform 1 0 12236 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_133
timestamp 1666464484
transform 1 0 13340 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1666464484
transform 1 0 14444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_151
timestamp 1666464484
transform 1 0 14996 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_163
timestamp 1666464484
transform 1 0 16100 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_175
timestamp 1666464484
transform 1 0 17204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_179
timestamp 1666464484
transform 1 0 17572 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_209
timestamp 1666464484
transform 1 0 20332 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_211
timestamp 1666464484
transform 1 0 20516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_235
timestamp 1666464484
transform 1 0 22724 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_239
timestamp 1666464484
transform 1 0 23092 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_241
timestamp 1666464484
transform 1 0 23276 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_253
timestamp 1666464484
transform 1 0 24380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_265
timestamp 1666464484
transform 1 0 25484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_269
timestamp 1666464484
transform 1 0 25852 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_271
timestamp 1666464484
transform 1 0 26036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_283
timestamp 1666464484
transform 1 0 27140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_295
timestamp 1666464484
transform 1 0 28244 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_299
timestamp 1666464484
transform 1 0 28612 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_301
timestamp 1666464484
transform 1 0 28796 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_313
timestamp 1666464484
transform 1 0 29900 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_325
timestamp 1666464484
transform 1 0 31004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_329
timestamp 1666464484
transform 1 0 31372 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_331
timestamp 1666464484
transform 1 0 31556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_343
timestamp 1666464484
transform 1 0 32660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_355
timestamp 1666464484
transform 1 0 33764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_359
timestamp 1666464484
transform 1 0 34132 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1666464484
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1666464484
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_385
timestamp 1666464484
transform 1 0 36524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_389
timestamp 1666464484
transform 1 0 36892 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_391
timestamp 1666464484
transform 1 0 37076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_403
timestamp 1666464484
transform 1 0 38180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_415
timestamp 1666464484
transform 1 0 39284 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_419
timestamp 1666464484
transform 1 0 39652 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_421
timestamp 1666464484
transform 1 0 39836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_433
timestamp 1666464484
transform 1 0 40940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_445
timestamp 1666464484
transform 1 0 42044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_449
timestamp 1666464484
transform 1 0 42412 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_451
timestamp 1666464484
transform 1 0 42596 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_463
timestamp 1666464484
transform 1 0 43700 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_475
timestamp 1666464484
transform 1 0 44804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_479
timestamp 1666464484
transform 1 0 45172 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_481
timestamp 1666464484
transform 1 0 45356 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_493
timestamp 1666464484
transform 1 0 46460 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_505
timestamp 1666464484
transform 1 0 47564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_509
timestamp 1666464484
transform 1 0 47932 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_511
timestamp 1666464484
transform 1 0 48116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_523
timestamp 1666464484
transform 1 0 49220 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_535
timestamp 1666464484
transform 1 0 50324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_539
timestamp 1666464484
transform 1 0 50692 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1666464484
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_553
timestamp 1666464484
transform 1 0 51980 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_565
timestamp 1666464484
transform 1 0 53084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_569
timestamp 1666464484
transform 1 0 53452 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_571
timestamp 1666464484
transform 1 0 53636 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_583
timestamp 1666464484
transform 1 0 54740 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_595
timestamp 1666464484
transform 1 0 55844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_599
timestamp 1666464484
transform 1 0 56212 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_601
timestamp 1666464484
transform 1 0 56396 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_613
timestamp 1666464484
transform 1 0 57500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_16
timestamp 1666464484
transform 1 0 2576 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_28
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_40
timestamp 1666464484
transform 1 0 4784 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_44
timestamp 1666464484
transform 1 0 5152 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_46
timestamp 1666464484
transform 1 0 5336 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_58
timestamp 1666464484
transform 1 0 6440 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_70
timestamp 1666464484
transform 1 0 7544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_74
timestamp 1666464484
transform 1 0 7912 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_76
timestamp 1666464484
transform 1 0 8096 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_88
timestamp 1666464484
transform 1 0 9200 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_100
timestamp 1666464484
transform 1 0 10304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_104
timestamp 1666464484
transform 1 0 10672 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_106
timestamp 1666464484
transform 1 0 10856 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_118
timestamp 1666464484
transform 1 0 11960 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1666464484
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_134
timestamp 1666464484
transform 1 0 13432 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_136
timestamp 1666464484
transform 1 0 13616 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_148
timestamp 1666464484
transform 1 0 14720 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_160
timestamp 1666464484
transform 1 0 15824 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_164
timestamp 1666464484
transform 1 0 16192 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_166
timestamp 1666464484
transform 1 0 16376 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_178
timestamp 1666464484
transform 1 0 17480 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_190
timestamp 1666464484
transform 1 0 18584 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_194
timestamp 1666464484
transform 1 0 18952 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_196
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_208
timestamp 1666464484
transform 1 0 20240 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_220
timestamp 1666464484
transform 1 0 21344 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_224
timestamp 1666464484
transform 1 0 21712 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_226
timestamp 1666464484
transform 1 0 21896 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_238
timestamp 1666464484
transform 1 0 23000 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_250
timestamp 1666464484
transform 1 0 24104 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_254
timestamp 1666464484
transform 1 0 24472 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_256
timestamp 1666464484
transform 1 0 24656 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_268
timestamp 1666464484
transform 1 0 25760 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_280
timestamp 1666464484
transform 1 0 26864 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_284
timestamp 1666464484
transform 1 0 27232 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_286
timestamp 1666464484
transform 1 0 27416 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_298
timestamp 1666464484
transform 1 0 28520 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_310
timestamp 1666464484
transform 1 0 29624 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_314
timestamp 1666464484
transform 1 0 29992 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_316
timestamp 1666464484
transform 1 0 30176 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_328
timestamp 1666464484
transform 1 0 31280 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_340
timestamp 1666464484
transform 1 0 32384 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_344
timestamp 1666464484
transform 1 0 32752 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_346
timestamp 1666464484
transform 1 0 32936 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_358
timestamp 1666464484
transform 1 0 34040 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_370
timestamp 1666464484
transform 1 0 35144 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_374
timestamp 1666464484
transform 1 0 35512 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_376
timestamp 1666464484
transform 1 0 35696 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_388
timestamp 1666464484
transform 1 0 36800 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_400
timestamp 1666464484
transform 1 0 37904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_404
timestamp 1666464484
transform 1 0 38272 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_406
timestamp 1666464484
transform 1 0 38456 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_418
timestamp 1666464484
transform 1 0 39560 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_430
timestamp 1666464484
transform 1 0 40664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_434
timestamp 1666464484
transform 1 0 41032 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_436
timestamp 1666464484
transform 1 0 41216 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_448
timestamp 1666464484
transform 1 0 42320 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_460
timestamp 1666464484
transform 1 0 43424 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_464
timestamp 1666464484
transform 1 0 43792 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_466
timestamp 1666464484
transform 1 0 43976 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_478
timestamp 1666464484
transform 1 0 45080 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_490
timestamp 1666464484
transform 1 0 46184 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_494
timestamp 1666464484
transform 1 0 46552 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_496
timestamp 1666464484
transform 1 0 46736 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_508
timestamp 1666464484
transform 1 0 47840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_520
timestamp 1666464484
transform 1 0 48944 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_524
timestamp 1666464484
transform 1 0 49312 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_526
timestamp 1666464484
transform 1 0 49496 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_538
timestamp 1666464484
transform 1 0 50600 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_550
timestamp 1666464484
transform 1 0 51704 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_554
timestamp 1666464484
transform 1 0 52072 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_556
timestamp 1666464484
transform 1 0 52256 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_568
timestamp 1666464484
transform 1 0 53360 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_580
timestamp 1666464484
transform 1 0 54464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_584
timestamp 1666464484
transform 1 0 54832 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_586
timestamp 1666464484
transform 1 0 55016 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_598
timestamp 1666464484
transform 1 0 56120 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_610
timestamp 1666464484
transform 1 0 57224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_614
timestamp 1666464484
transform 1 0 57592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_616
timestamp 1666464484
transform 1 0 57776 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_624
timestamp 1666464484
transform 1 0 58512 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_31
timestamp 1666464484
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_43
timestamp 1666464484
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_59
timestamp 1666464484
transform 1 0 6532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_61
timestamp 1666464484
transform 1 0 6716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_73
timestamp 1666464484
transform 1 0 7820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_85
timestamp 1666464484
transform 1 0 8924 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_89
timestamp 1666464484
transform 1 0 9292 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_91
timestamp 1666464484
transform 1 0 9476 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_103
timestamp 1666464484
transform 1 0 10580 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1666464484
transform 1 0 11684 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1666464484
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_121
timestamp 1666464484
transform 1 0 12236 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_133
timestamp 1666464484
transform 1 0 13340 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_145
timestamp 1666464484
transform 1 0 14444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_151
timestamp 1666464484
transform 1 0 14996 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_163
timestamp 1666464484
transform 1 0 16100 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_175
timestamp 1666464484
transform 1 0 17204 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_179
timestamp 1666464484
transform 1 0 17572 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_209
timestamp 1666464484
transform 1 0 20332 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_211
timestamp 1666464484
transform 1 0 20516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_235
timestamp 1666464484
transform 1 0 22724 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_239
timestamp 1666464484
transform 1 0 23092 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_241
timestamp 1666464484
transform 1 0 23276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_253
timestamp 1666464484
transform 1 0 24380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_265
timestamp 1666464484
transform 1 0 25484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_269
timestamp 1666464484
transform 1 0 25852 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_271
timestamp 1666464484
transform 1 0 26036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_283
timestamp 1666464484
transform 1 0 27140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_295
timestamp 1666464484
transform 1 0 28244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_299
timestamp 1666464484
transform 1 0 28612 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_301
timestamp 1666464484
transform 1 0 28796 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_313
timestamp 1666464484
transform 1 0 29900 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_325
timestamp 1666464484
transform 1 0 31004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_329
timestamp 1666464484
transform 1 0 31372 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_331
timestamp 1666464484
transform 1 0 31556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_343
timestamp 1666464484
transform 1 0 32660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_355
timestamp 1666464484
transform 1 0 33764 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_359
timestamp 1666464484
transform 1 0 34132 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1666464484
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1666464484
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_385
timestamp 1666464484
transform 1 0 36524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_389
timestamp 1666464484
transform 1 0 36892 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_391
timestamp 1666464484
transform 1 0 37076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_403
timestamp 1666464484
transform 1 0 38180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_415
timestamp 1666464484
transform 1 0 39284 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_419
timestamp 1666464484
transform 1 0 39652 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_421
timestamp 1666464484
transform 1 0 39836 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_433
timestamp 1666464484
transform 1 0 40940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_445
timestamp 1666464484
transform 1 0 42044 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_449
timestamp 1666464484
transform 1 0 42412 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_451
timestamp 1666464484
transform 1 0 42596 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_463
timestamp 1666464484
transform 1 0 43700 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_475
timestamp 1666464484
transform 1 0 44804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_479
timestamp 1666464484
transform 1 0 45172 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_481
timestamp 1666464484
transform 1 0 45356 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_493
timestamp 1666464484
transform 1 0 46460 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1666464484
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_509
timestamp 1666464484
transform 1 0 47932 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_511
timestamp 1666464484
transform 1 0 48116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_523
timestamp 1666464484
transform 1 0 49220 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_535
timestamp 1666464484
transform 1 0 50324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_539
timestamp 1666464484
transform 1 0 50692 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1666464484
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_553
timestamp 1666464484
transform 1 0 51980 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_565
timestamp 1666464484
transform 1 0 53084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_569
timestamp 1666464484
transform 1 0 53452 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_571
timestamp 1666464484
transform 1 0 53636 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_583
timestamp 1666464484
transform 1 0 54740 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_595
timestamp 1666464484
transform 1 0 55844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_599
timestamp 1666464484
transform 1 0 56212 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_601
timestamp 1666464484
transform 1 0 56396 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_613
timestamp 1666464484
transform 1 0 57500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_16
timestamp 1666464484
transform 1 0 2576 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_28
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_40
timestamp 1666464484
transform 1 0 4784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_44
timestamp 1666464484
transform 1 0 5152 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_46
timestamp 1666464484
transform 1 0 5336 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_58
timestamp 1666464484
transform 1 0 6440 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_70
timestamp 1666464484
transform 1 0 7544 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_74
timestamp 1666464484
transform 1 0 7912 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_76
timestamp 1666464484
transform 1 0 8096 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_88
timestamp 1666464484
transform 1 0 9200 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_100
timestamp 1666464484
transform 1 0 10304 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_104
timestamp 1666464484
transform 1 0 10672 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_106
timestamp 1666464484
transform 1 0 10856 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_118
timestamp 1666464484
transform 1 0 11960 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_130
timestamp 1666464484
transform 1 0 13064 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_134
timestamp 1666464484
transform 1 0 13432 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_136
timestamp 1666464484
transform 1 0 13616 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_148
timestamp 1666464484
transform 1 0 14720 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_160
timestamp 1666464484
transform 1 0 15824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_164
timestamp 1666464484
transform 1 0 16192 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_166
timestamp 1666464484
transform 1 0 16376 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_178
timestamp 1666464484
transform 1 0 17480 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_190
timestamp 1666464484
transform 1 0 18584 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_194
timestamp 1666464484
transform 1 0 18952 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_196
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_208
timestamp 1666464484
transform 1 0 20240 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_220
timestamp 1666464484
transform 1 0 21344 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_224
timestamp 1666464484
transform 1 0 21712 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_226
timestamp 1666464484
transform 1 0 21896 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_238
timestamp 1666464484
transform 1 0 23000 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_250
timestamp 1666464484
transform 1 0 24104 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_254
timestamp 1666464484
transform 1 0 24472 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_256
timestamp 1666464484
transform 1 0 24656 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_268
timestamp 1666464484
transform 1 0 25760 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_280
timestamp 1666464484
transform 1 0 26864 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_284
timestamp 1666464484
transform 1 0 27232 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_286
timestamp 1666464484
transform 1 0 27416 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_298
timestamp 1666464484
transform 1 0 28520 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_310
timestamp 1666464484
transform 1 0 29624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_314
timestamp 1666464484
transform 1 0 29992 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_316
timestamp 1666464484
transform 1 0 30176 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_328
timestamp 1666464484
transform 1 0 31280 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_340
timestamp 1666464484
transform 1 0 32384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_344
timestamp 1666464484
transform 1 0 32752 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_346
timestamp 1666464484
transform 1 0 32936 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_358
timestamp 1666464484
transform 1 0 34040 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_370
timestamp 1666464484
transform 1 0 35144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_374
timestamp 1666464484
transform 1 0 35512 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_376
timestamp 1666464484
transform 1 0 35696 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_388
timestamp 1666464484
transform 1 0 36800 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_400
timestamp 1666464484
transform 1 0 37904 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_404
timestamp 1666464484
transform 1 0 38272 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_406
timestamp 1666464484
transform 1 0 38456 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_418
timestamp 1666464484
transform 1 0 39560 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_430
timestamp 1666464484
transform 1 0 40664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_434
timestamp 1666464484
transform 1 0 41032 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_436
timestamp 1666464484
transform 1 0 41216 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_448
timestamp 1666464484
transform 1 0 42320 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_460
timestamp 1666464484
transform 1 0 43424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_464
timestamp 1666464484
transform 1 0 43792 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_466
timestamp 1666464484
transform 1 0 43976 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_478
timestamp 1666464484
transform 1 0 45080 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_490
timestamp 1666464484
transform 1 0 46184 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_494
timestamp 1666464484
transform 1 0 46552 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_496
timestamp 1666464484
transform 1 0 46736 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_508
timestamp 1666464484
transform 1 0 47840 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_520
timestamp 1666464484
transform 1 0 48944 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_524
timestamp 1666464484
transform 1 0 49312 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_526
timestamp 1666464484
transform 1 0 49496 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_538
timestamp 1666464484
transform 1 0 50600 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_550
timestamp 1666464484
transform 1 0 51704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_554
timestamp 1666464484
transform 1 0 52072 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_556
timestamp 1666464484
transform 1 0 52256 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_568
timestamp 1666464484
transform 1 0 53360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_580
timestamp 1666464484
transform 1 0 54464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_584
timestamp 1666464484
transform 1 0 54832 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_586
timestamp 1666464484
transform 1 0 55016 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_598
timestamp 1666464484
transform 1 0 56120 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_610
timestamp 1666464484
transform 1 0 57224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_614
timestamp 1666464484
transform 1 0 57592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_616
timestamp 1666464484
transform 1 0 57776 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_624
timestamp 1666464484
transform 1 0 58512 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_27
timestamp 1666464484
transform 1 0 3588 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_31
timestamp 1666464484
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_43
timestamp 1666464484
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_55
timestamp 1666464484
transform 1 0 6164 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_59
timestamp 1666464484
transform 1 0 6532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_61
timestamp 1666464484
transform 1 0 6716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_73
timestamp 1666464484
transform 1 0 7820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 1666464484
transform 1 0 8924 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_89
timestamp 1666464484
transform 1 0 9292 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_91
timestamp 1666464484
transform 1 0 9476 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_103
timestamp 1666464484
transform 1 0 10580 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1666464484
transform 1 0 11684 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_119
timestamp 1666464484
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_121
timestamp 1666464484
transform 1 0 12236 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_133
timestamp 1666464484
transform 1 0 13340 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_145
timestamp 1666464484
transform 1 0 14444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_151
timestamp 1666464484
transform 1 0 14996 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_163
timestamp 1666464484
transform 1 0 16100 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_175
timestamp 1666464484
transform 1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_179
timestamp 1666464484
transform 1 0 17572 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_209
timestamp 1666464484
transform 1 0 20332 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_211
timestamp 1666464484
transform 1 0 20516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_235
timestamp 1666464484
transform 1 0 22724 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_239
timestamp 1666464484
transform 1 0 23092 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_241
timestamp 1666464484
transform 1 0 23276 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_253
timestamp 1666464484
transform 1 0 24380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_265
timestamp 1666464484
transform 1 0 25484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_269
timestamp 1666464484
transform 1 0 25852 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_271
timestamp 1666464484
transform 1 0 26036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_283
timestamp 1666464484
transform 1 0 27140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_295
timestamp 1666464484
transform 1 0 28244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_299
timestamp 1666464484
transform 1 0 28612 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_301
timestamp 1666464484
transform 1 0 28796 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_313
timestamp 1666464484
transform 1 0 29900 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_325
timestamp 1666464484
transform 1 0 31004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_329
timestamp 1666464484
transform 1 0 31372 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_331
timestamp 1666464484
transform 1 0 31556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_343
timestamp 1666464484
transform 1 0 32660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_355
timestamp 1666464484
transform 1 0 33764 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_359
timestamp 1666464484
transform 1 0 34132 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1666464484
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1666464484
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_385
timestamp 1666464484
transform 1 0 36524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_389
timestamp 1666464484
transform 1 0 36892 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_391
timestamp 1666464484
transform 1 0 37076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_403
timestamp 1666464484
transform 1 0 38180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_415
timestamp 1666464484
transform 1 0 39284 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_419
timestamp 1666464484
transform 1 0 39652 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_421
timestamp 1666464484
transform 1 0 39836 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_433
timestamp 1666464484
transform 1 0 40940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_445
timestamp 1666464484
transform 1 0 42044 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_449
timestamp 1666464484
transform 1 0 42412 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_451
timestamp 1666464484
transform 1 0 42596 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_463
timestamp 1666464484
transform 1 0 43700 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_475
timestamp 1666464484
transform 1 0 44804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_479
timestamp 1666464484
transform 1 0 45172 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_481
timestamp 1666464484
transform 1 0 45356 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_493
timestamp 1666464484
transform 1 0 46460 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1666464484
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_509
timestamp 1666464484
transform 1 0 47932 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_511
timestamp 1666464484
transform 1 0 48116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_523
timestamp 1666464484
transform 1 0 49220 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_535
timestamp 1666464484
transform 1 0 50324 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_539
timestamp 1666464484
transform 1 0 50692 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1666464484
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_553
timestamp 1666464484
transform 1 0 51980 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_565
timestamp 1666464484
transform 1 0 53084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_569
timestamp 1666464484
transform 1 0 53452 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_571
timestamp 1666464484
transform 1 0 53636 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_583
timestamp 1666464484
transform 1 0 54740 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_595
timestamp 1666464484
transform 1 0 55844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_599
timestamp 1666464484
transform 1 0 56212 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_601
timestamp 1666464484
transform 1 0 56396 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_613
timestamp 1666464484
transform 1 0 57500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_16
timestamp 1666464484
transform 1 0 2576 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_28
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_40
timestamp 1666464484
transform 1 0 4784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_44
timestamp 1666464484
transform 1 0 5152 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_46
timestamp 1666464484
transform 1 0 5336 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_58
timestamp 1666464484
transform 1 0 6440 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_70
timestamp 1666464484
transform 1 0 7544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_74
timestamp 1666464484
transform 1 0 7912 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_76
timestamp 1666464484
transform 1 0 8096 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_88
timestamp 1666464484
transform 1 0 9200 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_100
timestamp 1666464484
transform 1 0 10304 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_104
timestamp 1666464484
transform 1 0 10672 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_106
timestamp 1666464484
transform 1 0 10856 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_118
timestamp 1666464484
transform 1 0 11960 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_130
timestamp 1666464484
transform 1 0 13064 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_134
timestamp 1666464484
transform 1 0 13432 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_136
timestamp 1666464484
transform 1 0 13616 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_148
timestamp 1666464484
transform 1 0 14720 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_160
timestamp 1666464484
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_164
timestamp 1666464484
transform 1 0 16192 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_166
timestamp 1666464484
transform 1 0 16376 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_178
timestamp 1666464484
transform 1 0 17480 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_190
timestamp 1666464484
transform 1 0 18584 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_194
timestamp 1666464484
transform 1 0 18952 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_196
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_208
timestamp 1666464484
transform 1 0 20240 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_220
timestamp 1666464484
transform 1 0 21344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_224
timestamp 1666464484
transform 1 0 21712 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_226
timestamp 1666464484
transform 1 0 21896 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_238
timestamp 1666464484
transform 1 0 23000 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_250
timestamp 1666464484
transform 1 0 24104 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_254
timestamp 1666464484
transform 1 0 24472 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_256
timestamp 1666464484
transform 1 0 24656 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_268
timestamp 1666464484
transform 1 0 25760 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_280
timestamp 1666464484
transform 1 0 26864 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_284
timestamp 1666464484
transform 1 0 27232 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_286
timestamp 1666464484
transform 1 0 27416 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_298
timestamp 1666464484
transform 1 0 28520 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_310
timestamp 1666464484
transform 1 0 29624 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_314
timestamp 1666464484
transform 1 0 29992 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_316
timestamp 1666464484
transform 1 0 30176 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_328
timestamp 1666464484
transform 1 0 31280 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_340
timestamp 1666464484
transform 1 0 32384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_344
timestamp 1666464484
transform 1 0 32752 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_346
timestamp 1666464484
transform 1 0 32936 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_358
timestamp 1666464484
transform 1 0 34040 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_370
timestamp 1666464484
transform 1 0 35144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_374
timestamp 1666464484
transform 1 0 35512 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_376
timestamp 1666464484
transform 1 0 35696 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_388
timestamp 1666464484
transform 1 0 36800 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_400
timestamp 1666464484
transform 1 0 37904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_404
timestamp 1666464484
transform 1 0 38272 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_406
timestamp 1666464484
transform 1 0 38456 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_418
timestamp 1666464484
transform 1 0 39560 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_430
timestamp 1666464484
transform 1 0 40664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_434
timestamp 1666464484
transform 1 0 41032 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_436
timestamp 1666464484
transform 1 0 41216 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_448
timestamp 1666464484
transform 1 0 42320 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_460
timestamp 1666464484
transform 1 0 43424 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_464
timestamp 1666464484
transform 1 0 43792 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_466
timestamp 1666464484
transform 1 0 43976 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_478
timestamp 1666464484
transform 1 0 45080 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_490
timestamp 1666464484
transform 1 0 46184 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_494
timestamp 1666464484
transform 1 0 46552 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_496
timestamp 1666464484
transform 1 0 46736 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_508
timestamp 1666464484
transform 1 0 47840 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_520
timestamp 1666464484
transform 1 0 48944 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_524
timestamp 1666464484
transform 1 0 49312 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_526
timestamp 1666464484
transform 1 0 49496 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_538
timestamp 1666464484
transform 1 0 50600 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_550
timestamp 1666464484
transform 1 0 51704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_554
timestamp 1666464484
transform 1 0 52072 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_556
timestamp 1666464484
transform 1 0 52256 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_568
timestamp 1666464484
transform 1 0 53360 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_580
timestamp 1666464484
transform 1 0 54464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_584
timestamp 1666464484
transform 1 0 54832 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_586
timestamp 1666464484
transform 1 0 55016 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_598
timestamp 1666464484
transform 1 0 56120 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_610
timestamp 1666464484
transform 1 0 57224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_614
timestamp 1666464484
transform 1 0 57592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_616
timestamp 1666464484
transform 1 0 57776 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_624
timestamp 1666464484
transform 1 0 58512 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_31
timestamp 1666464484
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_43
timestamp 1666464484
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_59
timestamp 1666464484
transform 1 0 6532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_61
timestamp 1666464484
transform 1 0 6716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_73
timestamp 1666464484
transform 1 0 7820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_85
timestamp 1666464484
transform 1 0 8924 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_89
timestamp 1666464484
transform 1 0 9292 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_91
timestamp 1666464484
transform 1 0 9476 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_103
timestamp 1666464484
transform 1 0 10580 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_115
timestamp 1666464484
transform 1 0 11684 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1666464484
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_121
timestamp 1666464484
transform 1 0 12236 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_133
timestamp 1666464484
transform 1 0 13340 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1666464484
transform 1 0 14444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_151
timestamp 1666464484
transform 1 0 14996 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_163
timestamp 1666464484
transform 1 0 16100 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_175
timestamp 1666464484
transform 1 0 17204 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_179
timestamp 1666464484
transform 1 0 17572 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_205
timestamp 1666464484
transform 1 0 19964 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_209
timestamp 1666464484
transform 1 0 20332 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_211
timestamp 1666464484
transform 1 0 20516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_235
timestamp 1666464484
transform 1 0 22724 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_239
timestamp 1666464484
transform 1 0 23092 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_241
timestamp 1666464484
transform 1 0 23276 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_253
timestamp 1666464484
transform 1 0 24380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_265
timestamp 1666464484
transform 1 0 25484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_269
timestamp 1666464484
transform 1 0 25852 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_271
timestamp 1666464484
transform 1 0 26036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_283
timestamp 1666464484
transform 1 0 27140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1666464484
transform 1 0 28244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_299
timestamp 1666464484
transform 1 0 28612 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_301
timestamp 1666464484
transform 1 0 28796 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_313
timestamp 1666464484
transform 1 0 29900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_325
timestamp 1666464484
transform 1 0 31004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_329
timestamp 1666464484
transform 1 0 31372 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_331
timestamp 1666464484
transform 1 0 31556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_343
timestamp 1666464484
transform 1 0 32660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_355
timestamp 1666464484
transform 1 0 33764 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_359
timestamp 1666464484
transform 1 0 34132 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1666464484
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1666464484
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_385
timestamp 1666464484
transform 1 0 36524 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_389
timestamp 1666464484
transform 1 0 36892 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_391
timestamp 1666464484
transform 1 0 37076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_403
timestamp 1666464484
transform 1 0 38180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_415
timestamp 1666464484
transform 1 0 39284 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_419
timestamp 1666464484
transform 1 0 39652 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_421
timestamp 1666464484
transform 1 0 39836 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_433
timestamp 1666464484
transform 1 0 40940 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_445
timestamp 1666464484
transform 1 0 42044 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_449
timestamp 1666464484
transform 1 0 42412 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_451
timestamp 1666464484
transform 1 0 42596 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_463
timestamp 1666464484
transform 1 0 43700 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_475
timestamp 1666464484
transform 1 0 44804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_479
timestamp 1666464484
transform 1 0 45172 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_481
timestamp 1666464484
transform 1 0 45356 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_493
timestamp 1666464484
transform 1 0 46460 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_505
timestamp 1666464484
transform 1 0 47564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_509
timestamp 1666464484
transform 1 0 47932 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_511
timestamp 1666464484
transform 1 0 48116 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_523
timestamp 1666464484
transform 1 0 49220 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_535
timestamp 1666464484
transform 1 0 50324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_539
timestamp 1666464484
transform 1 0 50692 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1666464484
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_553
timestamp 1666464484
transform 1 0 51980 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_565
timestamp 1666464484
transform 1 0 53084 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_569
timestamp 1666464484
transform 1 0 53452 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_571
timestamp 1666464484
transform 1 0 53636 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_583
timestamp 1666464484
transform 1 0 54740 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_595
timestamp 1666464484
transform 1 0 55844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_599
timestamp 1666464484
transform 1 0 56212 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_601
timestamp 1666464484
transform 1 0 56396 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_613
timestamp 1666464484
transform 1 0 57500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_16
timestamp 1666464484
transform 1 0 2576 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_28
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1666464484
transform 1 0 4784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_44
timestamp 1666464484
transform 1 0 5152 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_46
timestamp 1666464484
transform 1 0 5336 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_58
timestamp 1666464484
transform 1 0 6440 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_70
timestamp 1666464484
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_74
timestamp 1666464484
transform 1 0 7912 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_76
timestamp 1666464484
transform 1 0 8096 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_88
timestamp 1666464484
transform 1 0 9200 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_100
timestamp 1666464484
transform 1 0 10304 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_104
timestamp 1666464484
transform 1 0 10672 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_106
timestamp 1666464484
transform 1 0 10856 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_118
timestamp 1666464484
transform 1 0 11960 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_130
timestamp 1666464484
transform 1 0 13064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_134
timestamp 1666464484
transform 1 0 13432 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_136
timestamp 1666464484
transform 1 0 13616 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_148
timestamp 1666464484
transform 1 0 14720 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_160
timestamp 1666464484
transform 1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_164
timestamp 1666464484
transform 1 0 16192 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_166
timestamp 1666464484
transform 1 0 16376 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_178
timestamp 1666464484
transform 1 0 17480 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_190
timestamp 1666464484
transform 1 0 18584 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_194
timestamp 1666464484
transform 1 0 18952 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_196
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_208
timestamp 1666464484
transform 1 0 20240 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_220
timestamp 1666464484
transform 1 0 21344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_224
timestamp 1666464484
transform 1 0 21712 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_226
timestamp 1666464484
transform 1 0 21896 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_238
timestamp 1666464484
transform 1 0 23000 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_250
timestamp 1666464484
transform 1 0 24104 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_254
timestamp 1666464484
transform 1 0 24472 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_256
timestamp 1666464484
transform 1 0 24656 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_268
timestamp 1666464484
transform 1 0 25760 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_280
timestamp 1666464484
transform 1 0 26864 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_284
timestamp 1666464484
transform 1 0 27232 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_286
timestamp 1666464484
transform 1 0 27416 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_298
timestamp 1666464484
transform 1 0 28520 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_310
timestamp 1666464484
transform 1 0 29624 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_314
timestamp 1666464484
transform 1 0 29992 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_316
timestamp 1666464484
transform 1 0 30176 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_328
timestamp 1666464484
transform 1 0 31280 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_340
timestamp 1666464484
transform 1 0 32384 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_344
timestamp 1666464484
transform 1 0 32752 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_346
timestamp 1666464484
transform 1 0 32936 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_358
timestamp 1666464484
transform 1 0 34040 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_370
timestamp 1666464484
transform 1 0 35144 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_374
timestamp 1666464484
transform 1 0 35512 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_376
timestamp 1666464484
transform 1 0 35696 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_388
timestamp 1666464484
transform 1 0 36800 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_400
timestamp 1666464484
transform 1 0 37904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_404
timestamp 1666464484
transform 1 0 38272 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_406
timestamp 1666464484
transform 1 0 38456 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_418
timestamp 1666464484
transform 1 0 39560 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_430
timestamp 1666464484
transform 1 0 40664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_434
timestamp 1666464484
transform 1 0 41032 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_436
timestamp 1666464484
transform 1 0 41216 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_448
timestamp 1666464484
transform 1 0 42320 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_460
timestamp 1666464484
transform 1 0 43424 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_464
timestamp 1666464484
transform 1 0 43792 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_466
timestamp 1666464484
transform 1 0 43976 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_478
timestamp 1666464484
transform 1 0 45080 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_490
timestamp 1666464484
transform 1 0 46184 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_494
timestamp 1666464484
transform 1 0 46552 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_496
timestamp 1666464484
transform 1 0 46736 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_508
timestamp 1666464484
transform 1 0 47840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_520
timestamp 1666464484
transform 1 0 48944 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_524
timestamp 1666464484
transform 1 0 49312 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_526
timestamp 1666464484
transform 1 0 49496 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_538
timestamp 1666464484
transform 1 0 50600 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_550
timestamp 1666464484
transform 1 0 51704 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_554
timestamp 1666464484
transform 1 0 52072 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_556
timestamp 1666464484
transform 1 0 52256 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_568
timestamp 1666464484
transform 1 0 53360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_580
timestamp 1666464484
transform 1 0 54464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_584
timestamp 1666464484
transform 1 0 54832 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_586
timestamp 1666464484
transform 1 0 55016 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_598
timestamp 1666464484
transform 1 0 56120 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_610
timestamp 1666464484
transform 1 0 57224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_614
timestamp 1666464484
transform 1 0 57592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_616
timestamp 1666464484
transform 1 0 57776 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_624
timestamp 1666464484
transform 1 0 58512 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_31
timestamp 1666464484
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_43
timestamp 1666464484
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_59
timestamp 1666464484
transform 1 0 6532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_61
timestamp 1666464484
transform 1 0 6716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_73
timestamp 1666464484
transform 1 0 7820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_85
timestamp 1666464484
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_89
timestamp 1666464484
transform 1 0 9292 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_91
timestamp 1666464484
transform 1 0 9476 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_103
timestamp 1666464484
transform 1 0 10580 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_115
timestamp 1666464484
transform 1 0 11684 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1666464484
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_121
timestamp 1666464484
transform 1 0 12236 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_133
timestamp 1666464484
transform 1 0 13340 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_145
timestamp 1666464484
transform 1 0 14444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_151
timestamp 1666464484
transform 1 0 14996 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_163
timestamp 1666464484
transform 1 0 16100 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_175
timestamp 1666464484
transform 1 0 17204 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_179
timestamp 1666464484
transform 1 0 17572 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_209
timestamp 1666464484
transform 1 0 20332 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_211
timestamp 1666464484
transform 1 0 20516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_235
timestamp 1666464484
transform 1 0 22724 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_239
timestamp 1666464484
transform 1 0 23092 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_241
timestamp 1666464484
transform 1 0 23276 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_253
timestamp 1666464484
transform 1 0 24380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_265
timestamp 1666464484
transform 1 0 25484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_269
timestamp 1666464484
transform 1 0 25852 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_271
timestamp 1666464484
transform 1 0 26036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_283
timestamp 1666464484
transform 1 0 27140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_295
timestamp 1666464484
transform 1 0 28244 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_299
timestamp 1666464484
transform 1 0 28612 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_301
timestamp 1666464484
transform 1 0 28796 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_313
timestamp 1666464484
transform 1 0 29900 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_325
timestamp 1666464484
transform 1 0 31004 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_329
timestamp 1666464484
transform 1 0 31372 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_331
timestamp 1666464484
transform 1 0 31556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_343
timestamp 1666464484
transform 1 0 32660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_355
timestamp 1666464484
transform 1 0 33764 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_359
timestamp 1666464484
transform 1 0 34132 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1666464484
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1666464484
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_385
timestamp 1666464484
transform 1 0 36524 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_389
timestamp 1666464484
transform 1 0 36892 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_391
timestamp 1666464484
transform 1 0 37076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_403
timestamp 1666464484
transform 1 0 38180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_415
timestamp 1666464484
transform 1 0 39284 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_419
timestamp 1666464484
transform 1 0 39652 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_421
timestamp 1666464484
transform 1 0 39836 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_433
timestamp 1666464484
transform 1 0 40940 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_445
timestamp 1666464484
transform 1 0 42044 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_449
timestamp 1666464484
transform 1 0 42412 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_451
timestamp 1666464484
transform 1 0 42596 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_463
timestamp 1666464484
transform 1 0 43700 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_475
timestamp 1666464484
transform 1 0 44804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_479
timestamp 1666464484
transform 1 0 45172 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_481
timestamp 1666464484
transform 1 0 45356 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_493
timestamp 1666464484
transform 1 0 46460 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_505
timestamp 1666464484
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_509
timestamp 1666464484
transform 1 0 47932 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_511
timestamp 1666464484
transform 1 0 48116 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_523
timestamp 1666464484
transform 1 0 49220 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_535
timestamp 1666464484
transform 1 0 50324 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_539
timestamp 1666464484
transform 1 0 50692 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1666464484
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_553
timestamp 1666464484
transform 1 0 51980 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_565
timestamp 1666464484
transform 1 0 53084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_569
timestamp 1666464484
transform 1 0 53452 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_571
timestamp 1666464484
transform 1 0 53636 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_583
timestamp 1666464484
transform 1 0 54740 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_595
timestamp 1666464484
transform 1 0 55844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_599
timestamp 1666464484
transform 1 0 56212 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_601
timestamp 1666464484
transform 1 0 56396 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_613
timestamp 1666464484
transform 1 0 57500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_16
timestamp 1666464484
transform 1 0 2576 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_28
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_40
timestamp 1666464484
transform 1 0 4784 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_44
timestamp 1666464484
transform 1 0 5152 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_46
timestamp 1666464484
transform 1 0 5336 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_58
timestamp 1666464484
transform 1 0 6440 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_70
timestamp 1666464484
transform 1 0 7544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_74
timestamp 1666464484
transform 1 0 7912 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_76
timestamp 1666464484
transform 1 0 8096 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_88
timestamp 1666464484
transform 1 0 9200 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_100
timestamp 1666464484
transform 1 0 10304 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_104
timestamp 1666464484
transform 1 0 10672 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_106
timestamp 1666464484
transform 1 0 10856 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_118
timestamp 1666464484
transform 1 0 11960 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_130
timestamp 1666464484
transform 1 0 13064 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_134
timestamp 1666464484
transform 1 0 13432 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_136
timestamp 1666464484
transform 1 0 13616 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_148
timestamp 1666464484
transform 1 0 14720 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_160
timestamp 1666464484
transform 1 0 15824 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_164
timestamp 1666464484
transform 1 0 16192 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_166
timestamp 1666464484
transform 1 0 16376 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_178
timestamp 1666464484
transform 1 0 17480 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_190
timestamp 1666464484
transform 1 0 18584 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_194
timestamp 1666464484
transform 1 0 18952 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_196
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_208
timestamp 1666464484
transform 1 0 20240 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_220
timestamp 1666464484
transform 1 0 21344 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_224
timestamp 1666464484
transform 1 0 21712 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_226
timestamp 1666464484
transform 1 0 21896 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_238
timestamp 1666464484
transform 1 0 23000 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_250
timestamp 1666464484
transform 1 0 24104 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_254
timestamp 1666464484
transform 1 0 24472 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_256
timestamp 1666464484
transform 1 0 24656 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_268
timestamp 1666464484
transform 1 0 25760 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_280
timestamp 1666464484
transform 1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_284
timestamp 1666464484
transform 1 0 27232 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_286
timestamp 1666464484
transform 1 0 27416 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_298
timestamp 1666464484
transform 1 0 28520 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_310
timestamp 1666464484
transform 1 0 29624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_314
timestamp 1666464484
transform 1 0 29992 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_316
timestamp 1666464484
transform 1 0 30176 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_328
timestamp 1666464484
transform 1 0 31280 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_340
timestamp 1666464484
transform 1 0 32384 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_344
timestamp 1666464484
transform 1 0 32752 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_346
timestamp 1666464484
transform 1 0 32936 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_358
timestamp 1666464484
transform 1 0 34040 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_370
timestamp 1666464484
transform 1 0 35144 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_374
timestamp 1666464484
transform 1 0 35512 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_376
timestamp 1666464484
transform 1 0 35696 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_388
timestamp 1666464484
transform 1 0 36800 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_400
timestamp 1666464484
transform 1 0 37904 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_404
timestamp 1666464484
transform 1 0 38272 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_406
timestamp 1666464484
transform 1 0 38456 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_418
timestamp 1666464484
transform 1 0 39560 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_430
timestamp 1666464484
transform 1 0 40664 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_434
timestamp 1666464484
transform 1 0 41032 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_436
timestamp 1666464484
transform 1 0 41216 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_448
timestamp 1666464484
transform 1 0 42320 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_460
timestamp 1666464484
transform 1 0 43424 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_464
timestamp 1666464484
transform 1 0 43792 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_466
timestamp 1666464484
transform 1 0 43976 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_478
timestamp 1666464484
transform 1 0 45080 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_490
timestamp 1666464484
transform 1 0 46184 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_494
timestamp 1666464484
transform 1 0 46552 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_496
timestamp 1666464484
transform 1 0 46736 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_508
timestamp 1666464484
transform 1 0 47840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_520
timestamp 1666464484
transform 1 0 48944 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_524
timestamp 1666464484
transform 1 0 49312 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_526
timestamp 1666464484
transform 1 0 49496 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_538
timestamp 1666464484
transform 1 0 50600 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_550
timestamp 1666464484
transform 1 0 51704 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_554
timestamp 1666464484
transform 1 0 52072 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_556
timestamp 1666464484
transform 1 0 52256 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_568
timestamp 1666464484
transform 1 0 53360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_580
timestamp 1666464484
transform 1 0 54464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_584
timestamp 1666464484
transform 1 0 54832 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_586
timestamp 1666464484
transform 1 0 55016 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_598
timestamp 1666464484
transform 1 0 56120 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_610
timestamp 1666464484
transform 1 0 57224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_614
timestamp 1666464484
transform 1 0 57592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_616
timestamp 1666464484
transform 1 0 57776 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_624
timestamp 1666464484
transform 1 0 58512 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_31
timestamp 1666464484
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_43
timestamp 1666464484
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_59
timestamp 1666464484
transform 1 0 6532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_61
timestamp 1666464484
transform 1 0 6716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_73
timestamp 1666464484
transform 1 0 7820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_85
timestamp 1666464484
transform 1 0 8924 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1666464484
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_91
timestamp 1666464484
transform 1 0 9476 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_103
timestamp 1666464484
transform 1 0 10580 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_115
timestamp 1666464484
transform 1 0 11684 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 1666464484
transform 1 0 12052 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_121
timestamp 1666464484
transform 1 0 12236 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_133
timestamp 1666464484
transform 1 0 13340 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_145
timestamp 1666464484
transform 1 0 14444 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_151
timestamp 1666464484
transform 1 0 14996 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_163
timestamp 1666464484
transform 1 0 16100 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_175
timestamp 1666464484
transform 1 0 17204 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_179
timestamp 1666464484
transform 1 0 17572 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_205
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_209
timestamp 1666464484
transform 1 0 20332 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_211
timestamp 1666464484
transform 1 0 20516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_235
timestamp 1666464484
transform 1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_239
timestamp 1666464484
transform 1 0 23092 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_241
timestamp 1666464484
transform 1 0 23276 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_253
timestamp 1666464484
transform 1 0 24380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_265
timestamp 1666464484
transform 1 0 25484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_269
timestamp 1666464484
transform 1 0 25852 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_271
timestamp 1666464484
transform 1 0 26036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_283
timestamp 1666464484
transform 1 0 27140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_295
timestamp 1666464484
transform 1 0 28244 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_299
timestamp 1666464484
transform 1 0 28612 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_301
timestamp 1666464484
transform 1 0 28796 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_313
timestamp 1666464484
transform 1 0 29900 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_325
timestamp 1666464484
transform 1 0 31004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_329
timestamp 1666464484
transform 1 0 31372 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_331
timestamp 1666464484
transform 1 0 31556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_343
timestamp 1666464484
transform 1 0 32660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_355
timestamp 1666464484
transform 1 0 33764 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_359
timestamp 1666464484
transform 1 0 34132 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1666464484
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1666464484
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_385
timestamp 1666464484
transform 1 0 36524 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_389
timestamp 1666464484
transform 1 0 36892 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_391
timestamp 1666464484
transform 1 0 37076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_403
timestamp 1666464484
transform 1 0 38180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_415
timestamp 1666464484
transform 1 0 39284 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_419
timestamp 1666464484
transform 1 0 39652 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_421
timestamp 1666464484
transform 1 0 39836 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_433
timestamp 1666464484
transform 1 0 40940 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_445
timestamp 1666464484
transform 1 0 42044 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_449
timestamp 1666464484
transform 1 0 42412 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_451
timestamp 1666464484
transform 1 0 42596 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_463
timestamp 1666464484
transform 1 0 43700 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_475
timestamp 1666464484
transform 1 0 44804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_479
timestamp 1666464484
transform 1 0 45172 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_481
timestamp 1666464484
transform 1 0 45356 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_493
timestamp 1666464484
transform 1 0 46460 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_505
timestamp 1666464484
transform 1 0 47564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_509
timestamp 1666464484
transform 1 0 47932 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_511
timestamp 1666464484
transform 1 0 48116 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_523
timestamp 1666464484
transform 1 0 49220 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_535
timestamp 1666464484
transform 1 0 50324 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_539
timestamp 1666464484
transform 1 0 50692 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1666464484
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_553
timestamp 1666464484
transform 1 0 51980 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_565
timestamp 1666464484
transform 1 0 53084 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_569
timestamp 1666464484
transform 1 0 53452 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_571
timestamp 1666464484
transform 1 0 53636 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_583
timestamp 1666464484
transform 1 0 54740 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_595
timestamp 1666464484
transform 1 0 55844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_599
timestamp 1666464484
transform 1 0 56212 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_601
timestamp 1666464484
transform 1 0 56396 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_613
timestamp 1666464484
transform 1 0 57500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_16
timestamp 1666464484
transform 1 0 2576 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_28
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_40
timestamp 1666464484
transform 1 0 4784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_44
timestamp 1666464484
transform 1 0 5152 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_46
timestamp 1666464484
transform 1 0 5336 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_58
timestamp 1666464484
transform 1 0 6440 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_70
timestamp 1666464484
transform 1 0 7544 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_74
timestamp 1666464484
transform 1 0 7912 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_76
timestamp 1666464484
transform 1 0 8096 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_88
timestamp 1666464484
transform 1 0 9200 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_100
timestamp 1666464484
transform 1 0 10304 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_104
timestamp 1666464484
transform 1 0 10672 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_106
timestamp 1666464484
transform 1 0 10856 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_118
timestamp 1666464484
transform 1 0 11960 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_130
timestamp 1666464484
transform 1 0 13064 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_134
timestamp 1666464484
transform 1 0 13432 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_136
timestamp 1666464484
transform 1 0 13616 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_148
timestamp 1666464484
transform 1 0 14720 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_160
timestamp 1666464484
transform 1 0 15824 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_164
timestamp 1666464484
transform 1 0 16192 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_166
timestamp 1666464484
transform 1 0 16376 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_178
timestamp 1666464484
transform 1 0 17480 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_190
timestamp 1666464484
transform 1 0 18584 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_194
timestamp 1666464484
transform 1 0 18952 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_196
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_208
timestamp 1666464484
transform 1 0 20240 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_220
timestamp 1666464484
transform 1 0 21344 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_224
timestamp 1666464484
transform 1 0 21712 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_226
timestamp 1666464484
transform 1 0 21896 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_238
timestamp 1666464484
transform 1 0 23000 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_250
timestamp 1666464484
transform 1 0 24104 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_254
timestamp 1666464484
transform 1 0 24472 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_256
timestamp 1666464484
transform 1 0 24656 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_268
timestamp 1666464484
transform 1 0 25760 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_280
timestamp 1666464484
transform 1 0 26864 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_284
timestamp 1666464484
transform 1 0 27232 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_286
timestamp 1666464484
transform 1 0 27416 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_298
timestamp 1666464484
transform 1 0 28520 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_310
timestamp 1666464484
transform 1 0 29624 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_314
timestamp 1666464484
transform 1 0 29992 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_316
timestamp 1666464484
transform 1 0 30176 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_328
timestamp 1666464484
transform 1 0 31280 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_340
timestamp 1666464484
transform 1 0 32384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_344
timestamp 1666464484
transform 1 0 32752 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_346
timestamp 1666464484
transform 1 0 32936 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_358
timestamp 1666464484
transform 1 0 34040 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_370
timestamp 1666464484
transform 1 0 35144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_374
timestamp 1666464484
transform 1 0 35512 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_376
timestamp 1666464484
transform 1 0 35696 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_388
timestamp 1666464484
transform 1 0 36800 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_400
timestamp 1666464484
transform 1 0 37904 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_404
timestamp 1666464484
transform 1 0 38272 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_406
timestamp 1666464484
transform 1 0 38456 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_418
timestamp 1666464484
transform 1 0 39560 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_430
timestamp 1666464484
transform 1 0 40664 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_434
timestamp 1666464484
transform 1 0 41032 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_436
timestamp 1666464484
transform 1 0 41216 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_448
timestamp 1666464484
transform 1 0 42320 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_460
timestamp 1666464484
transform 1 0 43424 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_464
timestamp 1666464484
transform 1 0 43792 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_466
timestamp 1666464484
transform 1 0 43976 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_478
timestamp 1666464484
transform 1 0 45080 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_490
timestamp 1666464484
transform 1 0 46184 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_494
timestamp 1666464484
transform 1 0 46552 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_496
timestamp 1666464484
transform 1 0 46736 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_508
timestamp 1666464484
transform 1 0 47840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_520
timestamp 1666464484
transform 1 0 48944 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_524
timestamp 1666464484
transform 1 0 49312 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_526
timestamp 1666464484
transform 1 0 49496 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_538
timestamp 1666464484
transform 1 0 50600 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_550
timestamp 1666464484
transform 1 0 51704 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_554
timestamp 1666464484
transform 1 0 52072 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_556
timestamp 1666464484
transform 1 0 52256 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_568
timestamp 1666464484
transform 1 0 53360 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_580
timestamp 1666464484
transform 1 0 54464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_584
timestamp 1666464484
transform 1 0 54832 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_586
timestamp 1666464484
transform 1 0 55016 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_598
timestamp 1666464484
transform 1 0 56120 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_610
timestamp 1666464484
transform 1 0 57224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_614
timestamp 1666464484
transform 1 0 57592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_616
timestamp 1666464484
transform 1 0 57776 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_624
timestamp 1666464484
transform 1 0 58512 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_31
timestamp 1666464484
transform 1 0 3956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_43
timestamp 1666464484
transform 1 0 5060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_55
timestamp 1666464484
transform 1 0 6164 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_59
timestamp 1666464484
transform 1 0 6532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_61
timestamp 1666464484
transform 1 0 6716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_73
timestamp 1666464484
transform 1 0 7820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_85
timestamp 1666464484
transform 1 0 8924 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_89
timestamp 1666464484
transform 1 0 9292 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_91
timestamp 1666464484
transform 1 0 9476 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_103
timestamp 1666464484
transform 1 0 10580 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_115
timestamp 1666464484
transform 1 0 11684 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1666464484
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_121
timestamp 1666464484
transform 1 0 12236 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_133
timestamp 1666464484
transform 1 0 13340 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_145
timestamp 1666464484
transform 1 0 14444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_151
timestamp 1666464484
transform 1 0 14996 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_163
timestamp 1666464484
transform 1 0 16100 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_175
timestamp 1666464484
transform 1 0 17204 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_179
timestamp 1666464484
transform 1 0 17572 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_209
timestamp 1666464484
transform 1 0 20332 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_211
timestamp 1666464484
transform 1 0 20516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_235
timestamp 1666464484
transform 1 0 22724 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_239
timestamp 1666464484
transform 1 0 23092 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_241
timestamp 1666464484
transform 1 0 23276 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_253
timestamp 1666464484
transform 1 0 24380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_265
timestamp 1666464484
transform 1 0 25484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_269
timestamp 1666464484
transform 1 0 25852 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_271
timestamp 1666464484
transform 1 0 26036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_283
timestamp 1666464484
transform 1 0 27140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_295
timestamp 1666464484
transform 1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_299
timestamp 1666464484
transform 1 0 28612 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_301
timestamp 1666464484
transform 1 0 28796 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_313
timestamp 1666464484
transform 1 0 29900 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_325
timestamp 1666464484
transform 1 0 31004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_329
timestamp 1666464484
transform 1 0 31372 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_331
timestamp 1666464484
transform 1 0 31556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_343
timestamp 1666464484
transform 1 0 32660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_355
timestamp 1666464484
transform 1 0 33764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_359
timestamp 1666464484
transform 1 0 34132 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1666464484
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1666464484
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_385
timestamp 1666464484
transform 1 0 36524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_389
timestamp 1666464484
transform 1 0 36892 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_391
timestamp 1666464484
transform 1 0 37076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_403
timestamp 1666464484
transform 1 0 38180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_415
timestamp 1666464484
transform 1 0 39284 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_419
timestamp 1666464484
transform 1 0 39652 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_421
timestamp 1666464484
transform 1 0 39836 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_433
timestamp 1666464484
transform 1 0 40940 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_445
timestamp 1666464484
transform 1 0 42044 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_449
timestamp 1666464484
transform 1 0 42412 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_451
timestamp 1666464484
transform 1 0 42596 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_463
timestamp 1666464484
transform 1 0 43700 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_475
timestamp 1666464484
transform 1 0 44804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_479
timestamp 1666464484
transform 1 0 45172 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_481
timestamp 1666464484
transform 1 0 45356 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_493
timestamp 1666464484
transform 1 0 46460 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_505
timestamp 1666464484
transform 1 0 47564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_509
timestamp 1666464484
transform 1 0 47932 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_511
timestamp 1666464484
transform 1 0 48116 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_523
timestamp 1666464484
transform 1 0 49220 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_535
timestamp 1666464484
transform 1 0 50324 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_539
timestamp 1666464484
transform 1 0 50692 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1666464484
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_553
timestamp 1666464484
transform 1 0 51980 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_565
timestamp 1666464484
transform 1 0 53084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_569
timestamp 1666464484
transform 1 0 53452 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_571
timestamp 1666464484
transform 1 0 53636 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_583
timestamp 1666464484
transform 1 0 54740 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_595
timestamp 1666464484
transform 1 0 55844 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_599
timestamp 1666464484
transform 1 0 56212 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_601
timestamp 1666464484
transform 1 0 56396 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_613
timestamp 1666464484
transform 1 0 57500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_16
timestamp 1666464484
transform 1 0 2576 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_28
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_40
timestamp 1666464484
transform 1 0 4784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_44
timestamp 1666464484
transform 1 0 5152 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_46
timestamp 1666464484
transform 1 0 5336 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_58
timestamp 1666464484
transform 1 0 6440 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_70
timestamp 1666464484
transform 1 0 7544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_74
timestamp 1666464484
transform 1 0 7912 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_76
timestamp 1666464484
transform 1 0 8096 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_88
timestamp 1666464484
transform 1 0 9200 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_100
timestamp 1666464484
transform 1 0 10304 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_104
timestamp 1666464484
transform 1 0 10672 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_106
timestamp 1666464484
transform 1 0 10856 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_118
timestamp 1666464484
transform 1 0 11960 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_130
timestamp 1666464484
transform 1 0 13064 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_134
timestamp 1666464484
transform 1 0 13432 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_136
timestamp 1666464484
transform 1 0 13616 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_148
timestamp 1666464484
transform 1 0 14720 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_160
timestamp 1666464484
transform 1 0 15824 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_164
timestamp 1666464484
transform 1 0 16192 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_166
timestamp 1666464484
transform 1 0 16376 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_178
timestamp 1666464484
transform 1 0 17480 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_190
timestamp 1666464484
transform 1 0 18584 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_194
timestamp 1666464484
transform 1 0 18952 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_196
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_208
timestamp 1666464484
transform 1 0 20240 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_220
timestamp 1666464484
transform 1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_224
timestamp 1666464484
transform 1 0 21712 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_226
timestamp 1666464484
transform 1 0 21896 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_238
timestamp 1666464484
transform 1 0 23000 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_250
timestamp 1666464484
transform 1 0 24104 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_254
timestamp 1666464484
transform 1 0 24472 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_256
timestamp 1666464484
transform 1 0 24656 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_268
timestamp 1666464484
transform 1 0 25760 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_280
timestamp 1666464484
transform 1 0 26864 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_284
timestamp 1666464484
transform 1 0 27232 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_286
timestamp 1666464484
transform 1 0 27416 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_298
timestamp 1666464484
transform 1 0 28520 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_310
timestamp 1666464484
transform 1 0 29624 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_314
timestamp 1666464484
transform 1 0 29992 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_316
timestamp 1666464484
transform 1 0 30176 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_328
timestamp 1666464484
transform 1 0 31280 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_340
timestamp 1666464484
transform 1 0 32384 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_344
timestamp 1666464484
transform 1 0 32752 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_346
timestamp 1666464484
transform 1 0 32936 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_358
timestamp 1666464484
transform 1 0 34040 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_370
timestamp 1666464484
transform 1 0 35144 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_374
timestamp 1666464484
transform 1 0 35512 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_376
timestamp 1666464484
transform 1 0 35696 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_388
timestamp 1666464484
transform 1 0 36800 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_400
timestamp 1666464484
transform 1 0 37904 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_404
timestamp 1666464484
transform 1 0 38272 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_406
timestamp 1666464484
transform 1 0 38456 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_418
timestamp 1666464484
transform 1 0 39560 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_430
timestamp 1666464484
transform 1 0 40664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_434
timestamp 1666464484
transform 1 0 41032 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_436
timestamp 1666464484
transform 1 0 41216 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_448
timestamp 1666464484
transform 1 0 42320 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_460
timestamp 1666464484
transform 1 0 43424 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_464
timestamp 1666464484
transform 1 0 43792 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_466
timestamp 1666464484
transform 1 0 43976 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_478
timestamp 1666464484
transform 1 0 45080 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_490
timestamp 1666464484
transform 1 0 46184 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_494
timestamp 1666464484
transform 1 0 46552 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_496
timestamp 1666464484
transform 1 0 46736 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_508
timestamp 1666464484
transform 1 0 47840 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_520
timestamp 1666464484
transform 1 0 48944 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_524
timestamp 1666464484
transform 1 0 49312 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_526
timestamp 1666464484
transform 1 0 49496 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_538
timestamp 1666464484
transform 1 0 50600 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_550
timestamp 1666464484
transform 1 0 51704 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_554
timestamp 1666464484
transform 1 0 52072 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_556
timestamp 1666464484
transform 1 0 52256 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_568
timestamp 1666464484
transform 1 0 53360 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_580
timestamp 1666464484
transform 1 0 54464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_584
timestamp 1666464484
transform 1 0 54832 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_586
timestamp 1666464484
transform 1 0 55016 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_598
timestamp 1666464484
transform 1 0 56120 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_610
timestamp 1666464484
transform 1 0 57224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_614
timestamp 1666464484
transform 1 0 57592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_616
timestamp 1666464484
transform 1 0 57776 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_624
timestamp 1666464484
transform 1 0 58512 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_31
timestamp 1666464484
transform 1 0 3956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_43
timestamp 1666464484
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_59
timestamp 1666464484
transform 1 0 6532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_61
timestamp 1666464484
transform 1 0 6716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_73
timestamp 1666464484
transform 1 0 7820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1666464484
transform 1 0 8924 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_89
timestamp 1666464484
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_91
timestamp 1666464484
transform 1 0 9476 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_103
timestamp 1666464484
transform 1 0 10580 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_115
timestamp 1666464484
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_119
timestamp 1666464484
transform 1 0 12052 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_121
timestamp 1666464484
transform 1 0 12236 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_133
timestamp 1666464484
transform 1 0 13340 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_145
timestamp 1666464484
transform 1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_151
timestamp 1666464484
transform 1 0 14996 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_163
timestamp 1666464484
transform 1 0 16100 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_175
timestamp 1666464484
transform 1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_179
timestamp 1666464484
transform 1 0 17572 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_205
timestamp 1666464484
transform 1 0 19964 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_209
timestamp 1666464484
transform 1 0 20332 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_211
timestamp 1666464484
transform 1 0 20516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_235
timestamp 1666464484
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_239
timestamp 1666464484
transform 1 0 23092 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_241
timestamp 1666464484
transform 1 0 23276 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_253
timestamp 1666464484
transform 1 0 24380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_265
timestamp 1666464484
transform 1 0 25484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_269
timestamp 1666464484
transform 1 0 25852 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_271
timestamp 1666464484
transform 1 0 26036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_283
timestamp 1666464484
transform 1 0 27140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_295
timestamp 1666464484
transform 1 0 28244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_299
timestamp 1666464484
transform 1 0 28612 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_301
timestamp 1666464484
transform 1 0 28796 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_313
timestamp 1666464484
transform 1 0 29900 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_325
timestamp 1666464484
transform 1 0 31004 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_329
timestamp 1666464484
transform 1 0 31372 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_331
timestamp 1666464484
transform 1 0 31556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_343
timestamp 1666464484
transform 1 0 32660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_355
timestamp 1666464484
transform 1 0 33764 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_359
timestamp 1666464484
transform 1 0 34132 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1666464484
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1666464484
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_385
timestamp 1666464484
transform 1 0 36524 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_389
timestamp 1666464484
transform 1 0 36892 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_391
timestamp 1666464484
transform 1 0 37076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_403
timestamp 1666464484
transform 1 0 38180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_415
timestamp 1666464484
transform 1 0 39284 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_419
timestamp 1666464484
transform 1 0 39652 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_421
timestamp 1666464484
transform 1 0 39836 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_433
timestamp 1666464484
transform 1 0 40940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_445
timestamp 1666464484
transform 1 0 42044 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_449
timestamp 1666464484
transform 1 0 42412 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_451
timestamp 1666464484
transform 1 0 42596 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_463
timestamp 1666464484
transform 1 0 43700 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_475
timestamp 1666464484
transform 1 0 44804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_479
timestamp 1666464484
transform 1 0 45172 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_481
timestamp 1666464484
transform 1 0 45356 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_493
timestamp 1666464484
transform 1 0 46460 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_505
timestamp 1666464484
transform 1 0 47564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_509
timestamp 1666464484
transform 1 0 47932 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_511
timestamp 1666464484
transform 1 0 48116 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_523
timestamp 1666464484
transform 1 0 49220 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_535
timestamp 1666464484
transform 1 0 50324 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_539
timestamp 1666464484
transform 1 0 50692 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1666464484
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_553
timestamp 1666464484
transform 1 0 51980 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_565
timestamp 1666464484
transform 1 0 53084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_569
timestamp 1666464484
transform 1 0 53452 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_571
timestamp 1666464484
transform 1 0 53636 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_583
timestamp 1666464484
transform 1 0 54740 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_595
timestamp 1666464484
transform 1 0 55844 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_599
timestamp 1666464484
transform 1 0 56212 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_601
timestamp 1666464484
transform 1 0 56396 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_613
timestamp 1666464484
transform 1 0 57500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_16
timestamp 1666464484
transform 1 0 2576 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_28
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1666464484
transform 1 0 4784 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_44
timestamp 1666464484
transform 1 0 5152 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_46
timestamp 1666464484
transform 1 0 5336 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_58
timestamp 1666464484
transform 1 0 6440 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_70
timestamp 1666464484
transform 1 0 7544 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_74
timestamp 1666464484
transform 1 0 7912 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_76
timestamp 1666464484
transform 1 0 8096 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_88
timestamp 1666464484
transform 1 0 9200 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_100
timestamp 1666464484
transform 1 0 10304 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_104
timestamp 1666464484
transform 1 0 10672 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_106
timestamp 1666464484
transform 1 0 10856 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_118
timestamp 1666464484
transform 1 0 11960 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_130
timestamp 1666464484
transform 1 0 13064 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_134
timestamp 1666464484
transform 1 0 13432 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_136
timestamp 1666464484
transform 1 0 13616 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_148
timestamp 1666464484
transform 1 0 14720 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_160
timestamp 1666464484
transform 1 0 15824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_164
timestamp 1666464484
transform 1 0 16192 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_166
timestamp 1666464484
transform 1 0 16376 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_178
timestamp 1666464484
transform 1 0 17480 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_190
timestamp 1666464484
transform 1 0 18584 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_194
timestamp 1666464484
transform 1 0 18952 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_196
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_208
timestamp 1666464484
transform 1 0 20240 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_220
timestamp 1666464484
transform 1 0 21344 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_224
timestamp 1666464484
transform 1 0 21712 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_226
timestamp 1666464484
transform 1 0 21896 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_238
timestamp 1666464484
transform 1 0 23000 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_250
timestamp 1666464484
transform 1 0 24104 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_254
timestamp 1666464484
transform 1 0 24472 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_256
timestamp 1666464484
transform 1 0 24656 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_268
timestamp 1666464484
transform 1 0 25760 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_280
timestamp 1666464484
transform 1 0 26864 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_284
timestamp 1666464484
transform 1 0 27232 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_286
timestamp 1666464484
transform 1 0 27416 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_298
timestamp 1666464484
transform 1 0 28520 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_310
timestamp 1666464484
transform 1 0 29624 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_314
timestamp 1666464484
transform 1 0 29992 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_316
timestamp 1666464484
transform 1 0 30176 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_328
timestamp 1666464484
transform 1 0 31280 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_340
timestamp 1666464484
transform 1 0 32384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_344
timestamp 1666464484
transform 1 0 32752 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_346
timestamp 1666464484
transform 1 0 32936 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_358
timestamp 1666464484
transform 1 0 34040 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_370
timestamp 1666464484
transform 1 0 35144 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_374
timestamp 1666464484
transform 1 0 35512 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_376
timestamp 1666464484
transform 1 0 35696 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_388
timestamp 1666464484
transform 1 0 36800 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_400
timestamp 1666464484
transform 1 0 37904 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_404
timestamp 1666464484
transform 1 0 38272 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_406
timestamp 1666464484
transform 1 0 38456 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_418
timestamp 1666464484
transform 1 0 39560 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_430
timestamp 1666464484
transform 1 0 40664 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_434
timestamp 1666464484
transform 1 0 41032 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_436
timestamp 1666464484
transform 1 0 41216 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_448
timestamp 1666464484
transform 1 0 42320 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_460
timestamp 1666464484
transform 1 0 43424 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_464
timestamp 1666464484
transform 1 0 43792 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_466
timestamp 1666464484
transform 1 0 43976 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_478
timestamp 1666464484
transform 1 0 45080 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_490
timestamp 1666464484
transform 1 0 46184 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_494
timestamp 1666464484
transform 1 0 46552 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_496
timestamp 1666464484
transform 1 0 46736 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_508
timestamp 1666464484
transform 1 0 47840 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_520
timestamp 1666464484
transform 1 0 48944 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_524
timestamp 1666464484
transform 1 0 49312 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_526
timestamp 1666464484
transform 1 0 49496 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_538
timestamp 1666464484
transform 1 0 50600 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_550
timestamp 1666464484
transform 1 0 51704 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_554
timestamp 1666464484
transform 1 0 52072 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_556
timestamp 1666464484
transform 1 0 52256 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_568
timestamp 1666464484
transform 1 0 53360 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_580
timestamp 1666464484
transform 1 0 54464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_584
timestamp 1666464484
transform 1 0 54832 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_586
timestamp 1666464484
transform 1 0 55016 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_598
timestamp 1666464484
transform 1 0 56120 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_610
timestamp 1666464484
transform 1 0 57224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_614
timestamp 1666464484
transform 1 0 57592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_616
timestamp 1666464484
transform 1 0 57776 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_624
timestamp 1666464484
transform 1 0 58512 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666464484
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_27
timestamp 1666464484
transform 1 0 3588 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_31
timestamp 1666464484
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1666464484
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_55
timestamp 1666464484
transform 1 0 6164 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_59
timestamp 1666464484
transform 1 0 6532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_61
timestamp 1666464484
transform 1 0 6716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_73
timestamp 1666464484
transform 1 0 7820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_85
timestamp 1666464484
transform 1 0 8924 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_89
timestamp 1666464484
transform 1 0 9292 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_91
timestamp 1666464484
transform 1 0 9476 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_103
timestamp 1666464484
transform 1 0 10580 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_115
timestamp 1666464484
transform 1 0 11684 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1666464484
transform 1 0 12052 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_121
timestamp 1666464484
transform 1 0 12236 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_133
timestamp 1666464484
transform 1 0 13340 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_145
timestamp 1666464484
transform 1 0 14444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_151
timestamp 1666464484
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_163
timestamp 1666464484
transform 1 0 16100 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_175
timestamp 1666464484
transform 1 0 17204 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_179
timestamp 1666464484
transform 1 0 17572 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_209
timestamp 1666464484
transform 1 0 20332 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_211
timestamp 1666464484
transform 1 0 20516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_235
timestamp 1666464484
transform 1 0 22724 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_239
timestamp 1666464484
transform 1 0 23092 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_241
timestamp 1666464484
transform 1 0 23276 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_253
timestamp 1666464484
transform 1 0 24380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_265
timestamp 1666464484
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_269
timestamp 1666464484
transform 1 0 25852 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_271
timestamp 1666464484
transform 1 0 26036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_283
timestamp 1666464484
transform 1 0 27140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_295
timestamp 1666464484
transform 1 0 28244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_299
timestamp 1666464484
transform 1 0 28612 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_301
timestamp 1666464484
transform 1 0 28796 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_313
timestamp 1666464484
transform 1 0 29900 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_325
timestamp 1666464484
transform 1 0 31004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_329
timestamp 1666464484
transform 1 0 31372 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_331
timestamp 1666464484
transform 1 0 31556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_343
timestamp 1666464484
transform 1 0 32660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_355
timestamp 1666464484
transform 1 0 33764 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_359
timestamp 1666464484
transform 1 0 34132 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1666464484
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1666464484
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_385
timestamp 1666464484
transform 1 0 36524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_389
timestamp 1666464484
transform 1 0 36892 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_391
timestamp 1666464484
transform 1 0 37076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_403
timestamp 1666464484
transform 1 0 38180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_415
timestamp 1666464484
transform 1 0 39284 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_419
timestamp 1666464484
transform 1 0 39652 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_421
timestamp 1666464484
transform 1 0 39836 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_433
timestamp 1666464484
transform 1 0 40940 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_445
timestamp 1666464484
transform 1 0 42044 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_449
timestamp 1666464484
transform 1 0 42412 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_451
timestamp 1666464484
transform 1 0 42596 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_463
timestamp 1666464484
transform 1 0 43700 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_475
timestamp 1666464484
transform 1 0 44804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_479
timestamp 1666464484
transform 1 0 45172 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_481
timestamp 1666464484
transform 1 0 45356 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_493
timestamp 1666464484
transform 1 0 46460 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_505
timestamp 1666464484
transform 1 0 47564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_509
timestamp 1666464484
transform 1 0 47932 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_511
timestamp 1666464484
transform 1 0 48116 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_523
timestamp 1666464484
transform 1 0 49220 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_535
timestamp 1666464484
transform 1 0 50324 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_539
timestamp 1666464484
transform 1 0 50692 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1666464484
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_553
timestamp 1666464484
transform 1 0 51980 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_565
timestamp 1666464484
transform 1 0 53084 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_569
timestamp 1666464484
transform 1 0 53452 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_571
timestamp 1666464484
transform 1 0 53636 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_583
timestamp 1666464484
transform 1 0 54740 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_595
timestamp 1666464484
transform 1 0 55844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_599
timestamp 1666464484
transform 1 0 56212 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_601
timestamp 1666464484
transform 1 0 56396 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_613
timestamp 1666464484
transform 1 0 57500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_16
timestamp 1666464484
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_28
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_40
timestamp 1666464484
transform 1 0 4784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_44
timestamp 1666464484
transform 1 0 5152 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_46
timestamp 1666464484
transform 1 0 5336 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_58
timestamp 1666464484
transform 1 0 6440 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_70
timestamp 1666464484
transform 1 0 7544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_74
timestamp 1666464484
transform 1 0 7912 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_76
timestamp 1666464484
transform 1 0 8096 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_88
timestamp 1666464484
transform 1 0 9200 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_100
timestamp 1666464484
transform 1 0 10304 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_104
timestamp 1666464484
transform 1 0 10672 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_106
timestamp 1666464484
transform 1 0 10856 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_118
timestamp 1666464484
transform 1 0 11960 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_130
timestamp 1666464484
transform 1 0 13064 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_134
timestamp 1666464484
transform 1 0 13432 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_136
timestamp 1666464484
transform 1 0 13616 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_148
timestamp 1666464484
transform 1 0 14720 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_160
timestamp 1666464484
transform 1 0 15824 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_164
timestamp 1666464484
transform 1 0 16192 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_166
timestamp 1666464484
transform 1 0 16376 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_178
timestamp 1666464484
transform 1 0 17480 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_190
timestamp 1666464484
transform 1 0 18584 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_194
timestamp 1666464484
transform 1 0 18952 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_196
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_208
timestamp 1666464484
transform 1 0 20240 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_220
timestamp 1666464484
transform 1 0 21344 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_224
timestamp 1666464484
transform 1 0 21712 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_226
timestamp 1666464484
transform 1 0 21896 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_238
timestamp 1666464484
transform 1 0 23000 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_250
timestamp 1666464484
transform 1 0 24104 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_254
timestamp 1666464484
transform 1 0 24472 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_256
timestamp 1666464484
transform 1 0 24656 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_268
timestamp 1666464484
transform 1 0 25760 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_280
timestamp 1666464484
transform 1 0 26864 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_284
timestamp 1666464484
transform 1 0 27232 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_286
timestamp 1666464484
transform 1 0 27416 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_298
timestamp 1666464484
transform 1 0 28520 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_310
timestamp 1666464484
transform 1 0 29624 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_314
timestamp 1666464484
transform 1 0 29992 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_316
timestamp 1666464484
transform 1 0 30176 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_328
timestamp 1666464484
transform 1 0 31280 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_340
timestamp 1666464484
transform 1 0 32384 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_344
timestamp 1666464484
transform 1 0 32752 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_346
timestamp 1666464484
transform 1 0 32936 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_358
timestamp 1666464484
transform 1 0 34040 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_370
timestamp 1666464484
transform 1 0 35144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_374
timestamp 1666464484
transform 1 0 35512 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_376
timestamp 1666464484
transform 1 0 35696 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_388
timestamp 1666464484
transform 1 0 36800 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_400
timestamp 1666464484
transform 1 0 37904 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_404
timestamp 1666464484
transform 1 0 38272 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_406
timestamp 1666464484
transform 1 0 38456 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_418
timestamp 1666464484
transform 1 0 39560 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_430
timestamp 1666464484
transform 1 0 40664 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_434
timestamp 1666464484
transform 1 0 41032 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_436
timestamp 1666464484
transform 1 0 41216 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_448
timestamp 1666464484
transform 1 0 42320 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_460
timestamp 1666464484
transform 1 0 43424 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_464
timestamp 1666464484
transform 1 0 43792 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_466
timestamp 1666464484
transform 1 0 43976 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_478
timestamp 1666464484
transform 1 0 45080 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_490
timestamp 1666464484
transform 1 0 46184 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_494
timestamp 1666464484
transform 1 0 46552 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_496
timestamp 1666464484
transform 1 0 46736 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_508
timestamp 1666464484
transform 1 0 47840 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_520
timestamp 1666464484
transform 1 0 48944 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_524
timestamp 1666464484
transform 1 0 49312 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_526
timestamp 1666464484
transform 1 0 49496 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_538
timestamp 1666464484
transform 1 0 50600 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_550
timestamp 1666464484
transform 1 0 51704 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_554
timestamp 1666464484
transform 1 0 52072 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_556
timestamp 1666464484
transform 1 0 52256 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_568
timestamp 1666464484
transform 1 0 53360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_580
timestamp 1666464484
transform 1 0 54464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_584
timestamp 1666464484
transform 1 0 54832 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_586
timestamp 1666464484
transform 1 0 55016 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_598
timestamp 1666464484
transform 1 0 56120 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_610
timestamp 1666464484
transform 1 0 57224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_614
timestamp 1666464484
transform 1 0 57592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_616
timestamp 1666464484
transform 1 0 57776 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_624
timestamp 1666464484
transform 1 0 58512 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_31
timestamp 1666464484
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_43
timestamp 1666464484
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_59
timestamp 1666464484
transform 1 0 6532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_61
timestamp 1666464484
transform 1 0 6716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_73
timestamp 1666464484
transform 1 0 7820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_85
timestamp 1666464484
transform 1 0 8924 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_89
timestamp 1666464484
transform 1 0 9292 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_91
timestamp 1666464484
transform 1 0 9476 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_103
timestamp 1666464484
transform 1 0 10580 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_115
timestamp 1666464484
transform 1 0 11684 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_119
timestamp 1666464484
transform 1 0 12052 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_121
timestamp 1666464484
transform 1 0 12236 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_133
timestamp 1666464484
transform 1 0 13340 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_145
timestamp 1666464484
transform 1 0 14444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_151
timestamp 1666464484
transform 1 0 14996 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_163
timestamp 1666464484
transform 1 0 16100 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_175
timestamp 1666464484
transform 1 0 17204 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_179
timestamp 1666464484
transform 1 0 17572 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_209
timestamp 1666464484
transform 1 0 20332 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_211
timestamp 1666464484
transform 1 0 20516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_235
timestamp 1666464484
transform 1 0 22724 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_239
timestamp 1666464484
transform 1 0 23092 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_241
timestamp 1666464484
transform 1 0 23276 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_253
timestamp 1666464484
transform 1 0 24380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_265
timestamp 1666464484
transform 1 0 25484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_269
timestamp 1666464484
transform 1 0 25852 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_271
timestamp 1666464484
transform 1 0 26036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_283
timestamp 1666464484
transform 1 0 27140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_295
timestamp 1666464484
transform 1 0 28244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_299
timestamp 1666464484
transform 1 0 28612 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_301
timestamp 1666464484
transform 1 0 28796 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_313
timestamp 1666464484
transform 1 0 29900 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_325
timestamp 1666464484
transform 1 0 31004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_329
timestamp 1666464484
transform 1 0 31372 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_331
timestamp 1666464484
transform 1 0 31556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_343
timestamp 1666464484
transform 1 0 32660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_355
timestamp 1666464484
transform 1 0 33764 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_359
timestamp 1666464484
transform 1 0 34132 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1666464484
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1666464484
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_385
timestamp 1666464484
transform 1 0 36524 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_389
timestamp 1666464484
transform 1 0 36892 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_391
timestamp 1666464484
transform 1 0 37076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_403
timestamp 1666464484
transform 1 0 38180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_415
timestamp 1666464484
transform 1 0 39284 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_419
timestamp 1666464484
transform 1 0 39652 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_421
timestamp 1666464484
transform 1 0 39836 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_433
timestamp 1666464484
transform 1 0 40940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_445
timestamp 1666464484
transform 1 0 42044 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_449
timestamp 1666464484
transform 1 0 42412 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_451
timestamp 1666464484
transform 1 0 42596 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_463
timestamp 1666464484
transform 1 0 43700 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_475
timestamp 1666464484
transform 1 0 44804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_479
timestamp 1666464484
transform 1 0 45172 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_481
timestamp 1666464484
transform 1 0 45356 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_493
timestamp 1666464484
transform 1 0 46460 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_505
timestamp 1666464484
transform 1 0 47564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_509
timestamp 1666464484
transform 1 0 47932 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_511
timestamp 1666464484
transform 1 0 48116 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_523
timestamp 1666464484
transform 1 0 49220 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_535
timestamp 1666464484
transform 1 0 50324 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_539
timestamp 1666464484
transform 1 0 50692 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1666464484
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_553
timestamp 1666464484
transform 1 0 51980 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_565
timestamp 1666464484
transform 1 0 53084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_569
timestamp 1666464484
transform 1 0 53452 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_571
timestamp 1666464484
transform 1 0 53636 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_583
timestamp 1666464484
transform 1 0 54740 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_595
timestamp 1666464484
transform 1 0 55844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_599
timestamp 1666464484
transform 1 0 56212 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_601
timestamp 1666464484
transform 1 0 56396 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_613
timestamp 1666464484
transform 1 0 57500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_16
timestamp 1666464484
transform 1 0 2576 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_28
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_40
timestamp 1666464484
transform 1 0 4784 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_44
timestamp 1666464484
transform 1 0 5152 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_46
timestamp 1666464484
transform 1 0 5336 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_58
timestamp 1666464484
transform 1 0 6440 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_70
timestamp 1666464484
transform 1 0 7544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_74
timestamp 1666464484
transform 1 0 7912 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_76
timestamp 1666464484
transform 1 0 8096 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_88
timestamp 1666464484
transform 1 0 9200 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_100
timestamp 1666464484
transform 1 0 10304 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_104
timestamp 1666464484
transform 1 0 10672 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_106
timestamp 1666464484
transform 1 0 10856 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_118
timestamp 1666464484
transform 1 0 11960 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_130
timestamp 1666464484
transform 1 0 13064 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_134
timestamp 1666464484
transform 1 0 13432 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_136
timestamp 1666464484
transform 1 0 13616 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_148
timestamp 1666464484
transform 1 0 14720 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_160
timestamp 1666464484
transform 1 0 15824 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_164
timestamp 1666464484
transform 1 0 16192 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_166
timestamp 1666464484
transform 1 0 16376 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_178
timestamp 1666464484
transform 1 0 17480 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_190
timestamp 1666464484
transform 1 0 18584 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_194
timestamp 1666464484
transform 1 0 18952 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_196
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_208
timestamp 1666464484
transform 1 0 20240 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_220
timestamp 1666464484
transform 1 0 21344 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_224
timestamp 1666464484
transform 1 0 21712 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_226
timestamp 1666464484
transform 1 0 21896 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_238
timestamp 1666464484
transform 1 0 23000 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_250
timestamp 1666464484
transform 1 0 24104 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_254
timestamp 1666464484
transform 1 0 24472 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_256
timestamp 1666464484
transform 1 0 24656 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_268
timestamp 1666464484
transform 1 0 25760 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_280
timestamp 1666464484
transform 1 0 26864 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_284
timestamp 1666464484
transform 1 0 27232 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_286
timestamp 1666464484
transform 1 0 27416 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_298
timestamp 1666464484
transform 1 0 28520 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_310
timestamp 1666464484
transform 1 0 29624 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_314
timestamp 1666464484
transform 1 0 29992 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_316
timestamp 1666464484
transform 1 0 30176 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_328
timestamp 1666464484
transform 1 0 31280 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_340
timestamp 1666464484
transform 1 0 32384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_344
timestamp 1666464484
transform 1 0 32752 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_346
timestamp 1666464484
transform 1 0 32936 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_358
timestamp 1666464484
transform 1 0 34040 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_370
timestamp 1666464484
transform 1 0 35144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_374
timestamp 1666464484
transform 1 0 35512 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_376
timestamp 1666464484
transform 1 0 35696 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_388
timestamp 1666464484
transform 1 0 36800 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_400
timestamp 1666464484
transform 1 0 37904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_404
timestamp 1666464484
transform 1 0 38272 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_406
timestamp 1666464484
transform 1 0 38456 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_418
timestamp 1666464484
transform 1 0 39560 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_430
timestamp 1666464484
transform 1 0 40664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_434
timestamp 1666464484
transform 1 0 41032 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_436
timestamp 1666464484
transform 1 0 41216 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_448
timestamp 1666464484
transform 1 0 42320 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_460
timestamp 1666464484
transform 1 0 43424 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_464
timestamp 1666464484
transform 1 0 43792 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_466
timestamp 1666464484
transform 1 0 43976 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_478
timestamp 1666464484
transform 1 0 45080 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_490
timestamp 1666464484
transform 1 0 46184 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_494
timestamp 1666464484
transform 1 0 46552 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_496
timestamp 1666464484
transform 1 0 46736 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_508
timestamp 1666464484
transform 1 0 47840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_520
timestamp 1666464484
transform 1 0 48944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_524
timestamp 1666464484
transform 1 0 49312 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_526
timestamp 1666464484
transform 1 0 49496 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_538
timestamp 1666464484
transform 1 0 50600 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_550
timestamp 1666464484
transform 1 0 51704 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_554
timestamp 1666464484
transform 1 0 52072 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_556
timestamp 1666464484
transform 1 0 52256 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_568
timestamp 1666464484
transform 1 0 53360 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_580
timestamp 1666464484
transform 1 0 54464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_584
timestamp 1666464484
transform 1 0 54832 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_586
timestamp 1666464484
transform 1 0 55016 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_598
timestamp 1666464484
transform 1 0 56120 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_610
timestamp 1666464484
transform 1 0 57224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_614
timestamp 1666464484
transform 1 0 57592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_616
timestamp 1666464484
transform 1 0 57776 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_624
timestamp 1666464484
transform 1 0 58512 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_31
timestamp 1666464484
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_43
timestamp 1666464484
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_59
timestamp 1666464484
transform 1 0 6532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_61
timestamp 1666464484
transform 1 0 6716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_73
timestamp 1666464484
transform 1 0 7820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_85
timestamp 1666464484
transform 1 0 8924 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_89
timestamp 1666464484
transform 1 0 9292 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_91
timestamp 1666464484
transform 1 0 9476 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_103
timestamp 1666464484
transform 1 0 10580 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_115
timestamp 1666464484
transform 1 0 11684 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1666464484
transform 1 0 12052 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_121
timestamp 1666464484
transform 1 0 12236 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_133
timestamp 1666464484
transform 1 0 13340 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_145
timestamp 1666464484
transform 1 0 14444 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_151
timestamp 1666464484
transform 1 0 14996 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_163
timestamp 1666464484
transform 1 0 16100 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_175
timestamp 1666464484
transform 1 0 17204 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_179
timestamp 1666464484
transform 1 0 17572 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1666464484
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_209
timestamp 1666464484
transform 1 0 20332 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_211
timestamp 1666464484
transform 1 0 20516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_235
timestamp 1666464484
transform 1 0 22724 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_239
timestamp 1666464484
transform 1 0 23092 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_241
timestamp 1666464484
transform 1 0 23276 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_253
timestamp 1666464484
transform 1 0 24380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_265
timestamp 1666464484
transform 1 0 25484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_269
timestamp 1666464484
transform 1 0 25852 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_271
timestamp 1666464484
transform 1 0 26036 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_283
timestamp 1666464484
transform 1 0 27140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_295
timestamp 1666464484
transform 1 0 28244 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_299
timestamp 1666464484
transform 1 0 28612 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_301
timestamp 1666464484
transform 1 0 28796 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_313
timestamp 1666464484
transform 1 0 29900 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_325
timestamp 1666464484
transform 1 0 31004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_329
timestamp 1666464484
transform 1 0 31372 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_331
timestamp 1666464484
transform 1 0 31556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_343
timestamp 1666464484
transform 1 0 32660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_355
timestamp 1666464484
transform 1 0 33764 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_359
timestamp 1666464484
transform 1 0 34132 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1666464484
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1666464484
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_385
timestamp 1666464484
transform 1 0 36524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_389
timestamp 1666464484
transform 1 0 36892 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_391
timestamp 1666464484
transform 1 0 37076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_403
timestamp 1666464484
transform 1 0 38180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_415
timestamp 1666464484
transform 1 0 39284 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_419
timestamp 1666464484
transform 1 0 39652 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_421
timestamp 1666464484
transform 1 0 39836 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_433
timestamp 1666464484
transform 1 0 40940 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_445
timestamp 1666464484
transform 1 0 42044 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_449
timestamp 1666464484
transform 1 0 42412 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_451
timestamp 1666464484
transform 1 0 42596 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_463
timestamp 1666464484
transform 1 0 43700 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_475
timestamp 1666464484
transform 1 0 44804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_479
timestamp 1666464484
transform 1 0 45172 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_481
timestamp 1666464484
transform 1 0 45356 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_493
timestamp 1666464484
transform 1 0 46460 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_505
timestamp 1666464484
transform 1 0 47564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_509
timestamp 1666464484
transform 1 0 47932 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_511
timestamp 1666464484
transform 1 0 48116 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_523
timestamp 1666464484
transform 1 0 49220 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_535
timestamp 1666464484
transform 1 0 50324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_539
timestamp 1666464484
transform 1 0 50692 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1666464484
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_553
timestamp 1666464484
transform 1 0 51980 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_565
timestamp 1666464484
transform 1 0 53084 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_569
timestamp 1666464484
transform 1 0 53452 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_571
timestamp 1666464484
transform 1 0 53636 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_583
timestamp 1666464484
transform 1 0 54740 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_595
timestamp 1666464484
transform 1 0 55844 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_599
timestamp 1666464484
transform 1 0 56212 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_601
timestamp 1666464484
transform 1 0 56396 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_613
timestamp 1666464484
transform 1 0 57500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_16
timestamp 1666464484
transform 1 0 2576 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_28
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_40
timestamp 1666464484
transform 1 0 4784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_44
timestamp 1666464484
transform 1 0 5152 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_46
timestamp 1666464484
transform 1 0 5336 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_58
timestamp 1666464484
transform 1 0 6440 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_70
timestamp 1666464484
transform 1 0 7544 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_74
timestamp 1666464484
transform 1 0 7912 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_76
timestamp 1666464484
transform 1 0 8096 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_88
timestamp 1666464484
transform 1 0 9200 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_100
timestamp 1666464484
transform 1 0 10304 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_104
timestamp 1666464484
transform 1 0 10672 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_106
timestamp 1666464484
transform 1 0 10856 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_118
timestamp 1666464484
transform 1 0 11960 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_130
timestamp 1666464484
transform 1 0 13064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_134
timestamp 1666464484
transform 1 0 13432 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_136
timestamp 1666464484
transform 1 0 13616 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_148
timestamp 1666464484
transform 1 0 14720 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_160
timestamp 1666464484
transform 1 0 15824 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_164
timestamp 1666464484
transform 1 0 16192 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_166
timestamp 1666464484
transform 1 0 16376 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_178
timestamp 1666464484
transform 1 0 17480 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_190
timestamp 1666464484
transform 1 0 18584 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_194
timestamp 1666464484
transform 1 0 18952 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_196
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_208
timestamp 1666464484
transform 1 0 20240 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_220
timestamp 1666464484
transform 1 0 21344 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_224
timestamp 1666464484
transform 1 0 21712 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_226
timestamp 1666464484
transform 1 0 21896 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_238
timestamp 1666464484
transform 1 0 23000 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_250
timestamp 1666464484
transform 1 0 24104 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_254
timestamp 1666464484
transform 1 0 24472 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_256
timestamp 1666464484
transform 1 0 24656 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_268
timestamp 1666464484
transform 1 0 25760 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_280
timestamp 1666464484
transform 1 0 26864 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_284
timestamp 1666464484
transform 1 0 27232 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_286
timestamp 1666464484
transform 1 0 27416 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_298
timestamp 1666464484
transform 1 0 28520 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_310
timestamp 1666464484
transform 1 0 29624 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_314
timestamp 1666464484
transform 1 0 29992 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_316
timestamp 1666464484
transform 1 0 30176 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_328
timestamp 1666464484
transform 1 0 31280 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_340
timestamp 1666464484
transform 1 0 32384 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_344
timestamp 1666464484
transform 1 0 32752 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_346
timestamp 1666464484
transform 1 0 32936 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_358
timestamp 1666464484
transform 1 0 34040 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_370
timestamp 1666464484
transform 1 0 35144 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_374
timestamp 1666464484
transform 1 0 35512 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_376
timestamp 1666464484
transform 1 0 35696 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_388
timestamp 1666464484
transform 1 0 36800 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_400
timestamp 1666464484
transform 1 0 37904 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_404
timestamp 1666464484
transform 1 0 38272 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_406
timestamp 1666464484
transform 1 0 38456 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_418
timestamp 1666464484
transform 1 0 39560 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_430
timestamp 1666464484
transform 1 0 40664 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_434
timestamp 1666464484
transform 1 0 41032 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_436
timestamp 1666464484
transform 1 0 41216 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_448
timestamp 1666464484
transform 1 0 42320 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_460
timestamp 1666464484
transform 1 0 43424 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_464
timestamp 1666464484
transform 1 0 43792 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_466
timestamp 1666464484
transform 1 0 43976 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_478
timestamp 1666464484
transform 1 0 45080 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_490
timestamp 1666464484
transform 1 0 46184 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_494
timestamp 1666464484
transform 1 0 46552 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_496
timestamp 1666464484
transform 1 0 46736 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_508
timestamp 1666464484
transform 1 0 47840 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_520
timestamp 1666464484
transform 1 0 48944 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_524
timestamp 1666464484
transform 1 0 49312 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_526
timestamp 1666464484
transform 1 0 49496 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_538
timestamp 1666464484
transform 1 0 50600 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_550
timestamp 1666464484
transform 1 0 51704 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_554
timestamp 1666464484
transform 1 0 52072 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_556
timestamp 1666464484
transform 1 0 52256 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_568
timestamp 1666464484
transform 1 0 53360 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_580
timestamp 1666464484
transform 1 0 54464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_584
timestamp 1666464484
transform 1 0 54832 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_586
timestamp 1666464484
transform 1 0 55016 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_598
timestamp 1666464484
transform 1 0 56120 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_610
timestamp 1666464484
transform 1 0 57224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_614
timestamp 1666464484
transform 1 0 57592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_616
timestamp 1666464484
transform 1 0 57776 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_624
timestamp 1666464484
transform 1 0 58512 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_27
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_31
timestamp 1666464484
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1666464484
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_55
timestamp 1666464484
transform 1 0 6164 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_59
timestamp 1666464484
transform 1 0 6532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_61
timestamp 1666464484
transform 1 0 6716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_73
timestamp 1666464484
transform 1 0 7820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_85
timestamp 1666464484
transform 1 0 8924 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_89
timestamp 1666464484
transform 1 0 9292 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_91
timestamp 1666464484
transform 1 0 9476 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_103
timestamp 1666464484
transform 1 0 10580 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_115
timestamp 1666464484
transform 1 0 11684 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 1666464484
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_121
timestamp 1666464484
transform 1 0 12236 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_133
timestamp 1666464484
transform 1 0 13340 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_145
timestamp 1666464484
transform 1 0 14444 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_151
timestamp 1666464484
transform 1 0 14996 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_163
timestamp 1666464484
transform 1 0 16100 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_175
timestamp 1666464484
transform 1 0 17204 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_179
timestamp 1666464484
transform 1 0 17572 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_205
timestamp 1666464484
transform 1 0 19964 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_209
timestamp 1666464484
transform 1 0 20332 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_211
timestamp 1666464484
transform 1 0 20516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_223
timestamp 1666464484
transform 1 0 21620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_235
timestamp 1666464484
transform 1 0 22724 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_239
timestamp 1666464484
transform 1 0 23092 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_241
timestamp 1666464484
transform 1 0 23276 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_253
timestamp 1666464484
transform 1 0 24380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_265
timestamp 1666464484
transform 1 0 25484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_269
timestamp 1666464484
transform 1 0 25852 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_271
timestamp 1666464484
transform 1 0 26036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_283
timestamp 1666464484
transform 1 0 27140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_295
timestamp 1666464484
transform 1 0 28244 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_299
timestamp 1666464484
transform 1 0 28612 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_301
timestamp 1666464484
transform 1 0 28796 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_313
timestamp 1666464484
transform 1 0 29900 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_325
timestamp 1666464484
transform 1 0 31004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_329
timestamp 1666464484
transform 1 0 31372 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_331
timestamp 1666464484
transform 1 0 31556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_343
timestamp 1666464484
transform 1 0 32660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_355
timestamp 1666464484
transform 1 0 33764 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_359
timestamp 1666464484
transform 1 0 34132 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1666464484
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1666464484
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_385
timestamp 1666464484
transform 1 0 36524 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_389
timestamp 1666464484
transform 1 0 36892 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_391
timestamp 1666464484
transform 1 0 37076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_403
timestamp 1666464484
transform 1 0 38180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_415
timestamp 1666464484
transform 1 0 39284 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_419
timestamp 1666464484
transform 1 0 39652 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_421
timestamp 1666464484
transform 1 0 39836 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_433
timestamp 1666464484
transform 1 0 40940 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_445
timestamp 1666464484
transform 1 0 42044 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_449
timestamp 1666464484
transform 1 0 42412 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_451
timestamp 1666464484
transform 1 0 42596 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_463
timestamp 1666464484
transform 1 0 43700 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_475
timestamp 1666464484
transform 1 0 44804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_479
timestamp 1666464484
transform 1 0 45172 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_481
timestamp 1666464484
transform 1 0 45356 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_493
timestamp 1666464484
transform 1 0 46460 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_505
timestamp 1666464484
transform 1 0 47564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_509
timestamp 1666464484
transform 1 0 47932 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_511
timestamp 1666464484
transform 1 0 48116 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_523
timestamp 1666464484
transform 1 0 49220 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_535
timestamp 1666464484
transform 1 0 50324 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_539
timestamp 1666464484
transform 1 0 50692 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1666464484
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_553
timestamp 1666464484
transform 1 0 51980 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_565
timestamp 1666464484
transform 1 0 53084 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_569
timestamp 1666464484
transform 1 0 53452 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_571
timestamp 1666464484
transform 1 0 53636 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_583
timestamp 1666464484
transform 1 0 54740 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_595
timestamp 1666464484
transform 1 0 55844 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_599
timestamp 1666464484
transform 1 0 56212 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_601
timestamp 1666464484
transform 1 0 56396 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_613
timestamp 1666464484
transform 1 0 57500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_16
timestamp 1666464484
transform 1 0 2576 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_28
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_40
timestamp 1666464484
transform 1 0 4784 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_44
timestamp 1666464484
transform 1 0 5152 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_46
timestamp 1666464484
transform 1 0 5336 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_58
timestamp 1666464484
transform 1 0 6440 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_70
timestamp 1666464484
transform 1 0 7544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_74
timestamp 1666464484
transform 1 0 7912 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_76
timestamp 1666464484
transform 1 0 8096 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_88
timestamp 1666464484
transform 1 0 9200 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_100
timestamp 1666464484
transform 1 0 10304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_104
timestamp 1666464484
transform 1 0 10672 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_106
timestamp 1666464484
transform 1 0 10856 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_118
timestamp 1666464484
transform 1 0 11960 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_130
timestamp 1666464484
transform 1 0 13064 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_134
timestamp 1666464484
transform 1 0 13432 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_136
timestamp 1666464484
transform 1 0 13616 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_148
timestamp 1666464484
transform 1 0 14720 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_160
timestamp 1666464484
transform 1 0 15824 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_164
timestamp 1666464484
transform 1 0 16192 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_166
timestamp 1666464484
transform 1 0 16376 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_178
timestamp 1666464484
transform 1 0 17480 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_190
timestamp 1666464484
transform 1 0 18584 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_194
timestamp 1666464484
transform 1 0 18952 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_196
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_208
timestamp 1666464484
transform 1 0 20240 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_220
timestamp 1666464484
transform 1 0 21344 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_224
timestamp 1666464484
transform 1 0 21712 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_226
timestamp 1666464484
transform 1 0 21896 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_238
timestamp 1666464484
transform 1 0 23000 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_250
timestamp 1666464484
transform 1 0 24104 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_254
timestamp 1666464484
transform 1 0 24472 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_256
timestamp 1666464484
transform 1 0 24656 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_268
timestamp 1666464484
transform 1 0 25760 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_280
timestamp 1666464484
transform 1 0 26864 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_284
timestamp 1666464484
transform 1 0 27232 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_286
timestamp 1666464484
transform 1 0 27416 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_298
timestamp 1666464484
transform 1 0 28520 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_310
timestamp 1666464484
transform 1 0 29624 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_314
timestamp 1666464484
transform 1 0 29992 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_316
timestamp 1666464484
transform 1 0 30176 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_328
timestamp 1666464484
transform 1 0 31280 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_340
timestamp 1666464484
transform 1 0 32384 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_344
timestamp 1666464484
transform 1 0 32752 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_346
timestamp 1666464484
transform 1 0 32936 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_358
timestamp 1666464484
transform 1 0 34040 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_370
timestamp 1666464484
transform 1 0 35144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_374
timestamp 1666464484
transform 1 0 35512 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_376
timestamp 1666464484
transform 1 0 35696 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_388
timestamp 1666464484
transform 1 0 36800 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_400
timestamp 1666464484
transform 1 0 37904 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_404
timestamp 1666464484
transform 1 0 38272 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_406
timestamp 1666464484
transform 1 0 38456 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_418
timestamp 1666464484
transform 1 0 39560 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_430
timestamp 1666464484
transform 1 0 40664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_434
timestamp 1666464484
transform 1 0 41032 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_436
timestamp 1666464484
transform 1 0 41216 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_448
timestamp 1666464484
transform 1 0 42320 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_460
timestamp 1666464484
transform 1 0 43424 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_464
timestamp 1666464484
transform 1 0 43792 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_466
timestamp 1666464484
transform 1 0 43976 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_478
timestamp 1666464484
transform 1 0 45080 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_490
timestamp 1666464484
transform 1 0 46184 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_494
timestamp 1666464484
transform 1 0 46552 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_496
timestamp 1666464484
transform 1 0 46736 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_508
timestamp 1666464484
transform 1 0 47840 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_520
timestamp 1666464484
transform 1 0 48944 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_524
timestamp 1666464484
transform 1 0 49312 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_526
timestamp 1666464484
transform 1 0 49496 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_538
timestamp 1666464484
transform 1 0 50600 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_550
timestamp 1666464484
transform 1 0 51704 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_554
timestamp 1666464484
transform 1 0 52072 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_556
timestamp 1666464484
transform 1 0 52256 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_568
timestamp 1666464484
transform 1 0 53360 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_580
timestamp 1666464484
transform 1 0 54464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_584
timestamp 1666464484
transform 1 0 54832 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_586
timestamp 1666464484
transform 1 0 55016 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_598
timestamp 1666464484
transform 1 0 56120 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_610
timestamp 1666464484
transform 1 0 57224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_614
timestamp 1666464484
transform 1 0 57592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_616
timestamp 1666464484
transform 1 0 57776 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_624
timestamp 1666464484
transform 1 0 58512 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666464484
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_27
timestamp 1666464484
transform 1 0 3588 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_31
timestamp 1666464484
transform 1 0 3956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_43
timestamp 1666464484
transform 1 0 5060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_55
timestamp 1666464484
transform 1 0 6164 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_59
timestamp 1666464484
transform 1 0 6532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_61
timestamp 1666464484
transform 1 0 6716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_73
timestamp 1666464484
transform 1 0 7820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_85
timestamp 1666464484
transform 1 0 8924 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_89
timestamp 1666464484
transform 1 0 9292 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_91
timestamp 1666464484
transform 1 0 9476 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_103
timestamp 1666464484
transform 1 0 10580 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_115
timestamp 1666464484
transform 1 0 11684 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_119
timestamp 1666464484
transform 1 0 12052 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_121
timestamp 1666464484
transform 1 0 12236 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_133
timestamp 1666464484
transform 1 0 13340 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_145
timestamp 1666464484
transform 1 0 14444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_151
timestamp 1666464484
transform 1 0 14996 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_163
timestamp 1666464484
transform 1 0 16100 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_175
timestamp 1666464484
transform 1 0 17204 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_179
timestamp 1666464484
transform 1 0 17572 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1666464484
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1666464484
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_205
timestamp 1666464484
transform 1 0 19964 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_209
timestamp 1666464484
transform 1 0 20332 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_211
timestamp 1666464484
transform 1 0 20516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_235
timestamp 1666464484
transform 1 0 22724 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_239
timestamp 1666464484
transform 1 0 23092 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_241
timestamp 1666464484
transform 1 0 23276 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_253
timestamp 1666464484
transform 1 0 24380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_265
timestamp 1666464484
transform 1 0 25484 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_269
timestamp 1666464484
transform 1 0 25852 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_271
timestamp 1666464484
transform 1 0 26036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_283
timestamp 1666464484
transform 1 0 27140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_295
timestamp 1666464484
transform 1 0 28244 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_299
timestamp 1666464484
transform 1 0 28612 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_301
timestamp 1666464484
transform 1 0 28796 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_313
timestamp 1666464484
transform 1 0 29900 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_325
timestamp 1666464484
transform 1 0 31004 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_329
timestamp 1666464484
transform 1 0 31372 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_331
timestamp 1666464484
transform 1 0 31556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_343
timestamp 1666464484
transform 1 0 32660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_355
timestamp 1666464484
transform 1 0 33764 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_359
timestamp 1666464484
transform 1 0 34132 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1666464484
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1666464484
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_385
timestamp 1666464484
transform 1 0 36524 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_389
timestamp 1666464484
transform 1 0 36892 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_391
timestamp 1666464484
transform 1 0 37076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_403
timestamp 1666464484
transform 1 0 38180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_415
timestamp 1666464484
transform 1 0 39284 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_419
timestamp 1666464484
transform 1 0 39652 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_421
timestamp 1666464484
transform 1 0 39836 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_433
timestamp 1666464484
transform 1 0 40940 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_445
timestamp 1666464484
transform 1 0 42044 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_449
timestamp 1666464484
transform 1 0 42412 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_451
timestamp 1666464484
transform 1 0 42596 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_463
timestamp 1666464484
transform 1 0 43700 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_475
timestamp 1666464484
transform 1 0 44804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_479
timestamp 1666464484
transform 1 0 45172 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_481
timestamp 1666464484
transform 1 0 45356 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_493
timestamp 1666464484
transform 1 0 46460 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_505
timestamp 1666464484
transform 1 0 47564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_509
timestamp 1666464484
transform 1 0 47932 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_511
timestamp 1666464484
transform 1 0 48116 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_523
timestamp 1666464484
transform 1 0 49220 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_535
timestamp 1666464484
transform 1 0 50324 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_539
timestamp 1666464484
transform 1 0 50692 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1666464484
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_553
timestamp 1666464484
transform 1 0 51980 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_565
timestamp 1666464484
transform 1 0 53084 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_569
timestamp 1666464484
transform 1 0 53452 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_571
timestamp 1666464484
transform 1 0 53636 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_583
timestamp 1666464484
transform 1 0 54740 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_595
timestamp 1666464484
transform 1 0 55844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_599
timestamp 1666464484
transform 1 0 56212 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_601
timestamp 1666464484
transform 1 0 56396 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_613
timestamp 1666464484
transform 1 0 57500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_16
timestamp 1666464484
transform 1 0 2576 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_28
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_40
timestamp 1666464484
transform 1 0 4784 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_44
timestamp 1666464484
transform 1 0 5152 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_46
timestamp 1666464484
transform 1 0 5336 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_58
timestamp 1666464484
transform 1 0 6440 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_70
timestamp 1666464484
transform 1 0 7544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_74
timestamp 1666464484
transform 1 0 7912 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_76
timestamp 1666464484
transform 1 0 8096 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_88
timestamp 1666464484
transform 1 0 9200 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_100
timestamp 1666464484
transform 1 0 10304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_104
timestamp 1666464484
transform 1 0 10672 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_106
timestamp 1666464484
transform 1 0 10856 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_118
timestamp 1666464484
transform 1 0 11960 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_130
timestamp 1666464484
transform 1 0 13064 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_134
timestamp 1666464484
transform 1 0 13432 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_136
timestamp 1666464484
transform 1 0 13616 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_148
timestamp 1666464484
transform 1 0 14720 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_160
timestamp 1666464484
transform 1 0 15824 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_164
timestamp 1666464484
transform 1 0 16192 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_166
timestamp 1666464484
transform 1 0 16376 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_178
timestamp 1666464484
transform 1 0 17480 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_190
timestamp 1666464484
transform 1 0 18584 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_194
timestamp 1666464484
transform 1 0 18952 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_196
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_208
timestamp 1666464484
transform 1 0 20240 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_220
timestamp 1666464484
transform 1 0 21344 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_224
timestamp 1666464484
transform 1 0 21712 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_226
timestamp 1666464484
transform 1 0 21896 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_238
timestamp 1666464484
transform 1 0 23000 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_250
timestamp 1666464484
transform 1 0 24104 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_254
timestamp 1666464484
transform 1 0 24472 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_256
timestamp 1666464484
transform 1 0 24656 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_268
timestamp 1666464484
transform 1 0 25760 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_280
timestamp 1666464484
transform 1 0 26864 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_284
timestamp 1666464484
transform 1 0 27232 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_286
timestamp 1666464484
transform 1 0 27416 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_298
timestamp 1666464484
transform 1 0 28520 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_310
timestamp 1666464484
transform 1 0 29624 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_314
timestamp 1666464484
transform 1 0 29992 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_316
timestamp 1666464484
transform 1 0 30176 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_328
timestamp 1666464484
transform 1 0 31280 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_340
timestamp 1666464484
transform 1 0 32384 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_344
timestamp 1666464484
transform 1 0 32752 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_346
timestamp 1666464484
transform 1 0 32936 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_358
timestamp 1666464484
transform 1 0 34040 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_370
timestamp 1666464484
transform 1 0 35144 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_374
timestamp 1666464484
transform 1 0 35512 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_376
timestamp 1666464484
transform 1 0 35696 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_388
timestamp 1666464484
transform 1 0 36800 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_400
timestamp 1666464484
transform 1 0 37904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_404
timestamp 1666464484
transform 1 0 38272 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_406
timestamp 1666464484
transform 1 0 38456 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_418
timestamp 1666464484
transform 1 0 39560 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_430
timestamp 1666464484
transform 1 0 40664 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_434
timestamp 1666464484
transform 1 0 41032 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_436
timestamp 1666464484
transform 1 0 41216 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_448
timestamp 1666464484
transform 1 0 42320 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_460
timestamp 1666464484
transform 1 0 43424 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_464
timestamp 1666464484
transform 1 0 43792 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_466
timestamp 1666464484
transform 1 0 43976 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_478
timestamp 1666464484
transform 1 0 45080 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_490
timestamp 1666464484
transform 1 0 46184 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_494
timestamp 1666464484
transform 1 0 46552 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_496
timestamp 1666464484
transform 1 0 46736 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_508
timestamp 1666464484
transform 1 0 47840 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_520
timestamp 1666464484
transform 1 0 48944 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_524
timestamp 1666464484
transform 1 0 49312 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_526
timestamp 1666464484
transform 1 0 49496 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_538
timestamp 1666464484
transform 1 0 50600 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_550
timestamp 1666464484
transform 1 0 51704 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_554
timestamp 1666464484
transform 1 0 52072 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_556
timestamp 1666464484
transform 1 0 52256 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_568
timestamp 1666464484
transform 1 0 53360 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_580
timestamp 1666464484
transform 1 0 54464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_584
timestamp 1666464484
transform 1 0 54832 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_586
timestamp 1666464484
transform 1 0 55016 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_598
timestamp 1666464484
transform 1 0 56120 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_610
timestamp 1666464484
transform 1 0 57224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_614
timestamp 1666464484
transform 1 0 57592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_616
timestamp 1666464484
transform 1 0 57776 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_624
timestamp 1666464484
transform 1 0 58512 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666464484
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_27
timestamp 1666464484
transform 1 0 3588 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_31
timestamp 1666464484
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_43
timestamp 1666464484
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_55
timestamp 1666464484
transform 1 0 6164 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_59
timestamp 1666464484
transform 1 0 6532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_61
timestamp 1666464484
transform 1 0 6716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_73
timestamp 1666464484
transform 1 0 7820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_85
timestamp 1666464484
transform 1 0 8924 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_89
timestamp 1666464484
transform 1 0 9292 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_91
timestamp 1666464484
transform 1 0 9476 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_103
timestamp 1666464484
transform 1 0 10580 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_115
timestamp 1666464484
transform 1 0 11684 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_119
timestamp 1666464484
transform 1 0 12052 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_121
timestamp 1666464484
transform 1 0 12236 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_133
timestamp 1666464484
transform 1 0 13340 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_145
timestamp 1666464484
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_151
timestamp 1666464484
transform 1 0 14996 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_163
timestamp 1666464484
transform 1 0 16100 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_175
timestamp 1666464484
transform 1 0 17204 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_179
timestamp 1666464484
transform 1 0 17572 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1666464484
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_205
timestamp 1666464484
transform 1 0 19964 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_209
timestamp 1666464484
transform 1 0 20332 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_211
timestamp 1666464484
transform 1 0 20516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_235
timestamp 1666464484
transform 1 0 22724 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_239
timestamp 1666464484
transform 1 0 23092 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_241
timestamp 1666464484
transform 1 0 23276 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_253
timestamp 1666464484
transform 1 0 24380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_265
timestamp 1666464484
transform 1 0 25484 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_269
timestamp 1666464484
transform 1 0 25852 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_271
timestamp 1666464484
transform 1 0 26036 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_283
timestamp 1666464484
transform 1 0 27140 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_295
timestamp 1666464484
transform 1 0 28244 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_299
timestamp 1666464484
transform 1 0 28612 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_301
timestamp 1666464484
transform 1 0 28796 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_313
timestamp 1666464484
transform 1 0 29900 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_325
timestamp 1666464484
transform 1 0 31004 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_329
timestamp 1666464484
transform 1 0 31372 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_331
timestamp 1666464484
transform 1 0 31556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_343
timestamp 1666464484
transform 1 0 32660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_355
timestamp 1666464484
transform 1 0 33764 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_359
timestamp 1666464484
transform 1 0 34132 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1666464484
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1666464484
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_385
timestamp 1666464484
transform 1 0 36524 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_389
timestamp 1666464484
transform 1 0 36892 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_391
timestamp 1666464484
transform 1 0 37076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_403
timestamp 1666464484
transform 1 0 38180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_415
timestamp 1666464484
transform 1 0 39284 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_419
timestamp 1666464484
transform 1 0 39652 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_421
timestamp 1666464484
transform 1 0 39836 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_433
timestamp 1666464484
transform 1 0 40940 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_445
timestamp 1666464484
transform 1 0 42044 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_449
timestamp 1666464484
transform 1 0 42412 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_451
timestamp 1666464484
transform 1 0 42596 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_463
timestamp 1666464484
transform 1 0 43700 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_475
timestamp 1666464484
transform 1 0 44804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_479
timestamp 1666464484
transform 1 0 45172 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_481
timestamp 1666464484
transform 1 0 45356 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_493
timestamp 1666464484
transform 1 0 46460 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_505
timestamp 1666464484
transform 1 0 47564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_509
timestamp 1666464484
transform 1 0 47932 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_511
timestamp 1666464484
transform 1 0 48116 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_523
timestamp 1666464484
transform 1 0 49220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_535
timestamp 1666464484
transform 1 0 50324 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_539
timestamp 1666464484
transform 1 0 50692 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1666464484
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_553
timestamp 1666464484
transform 1 0 51980 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_565
timestamp 1666464484
transform 1 0 53084 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_569
timestamp 1666464484
transform 1 0 53452 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_571
timestamp 1666464484
transform 1 0 53636 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_583
timestamp 1666464484
transform 1 0 54740 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_595
timestamp 1666464484
transform 1 0 55844 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_599
timestamp 1666464484
transform 1 0 56212 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_601
timestamp 1666464484
transform 1 0 56396 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_613
timestamp 1666464484
transform 1 0 57500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_16
timestamp 1666464484
transform 1 0 2576 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_28
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_40
timestamp 1666464484
transform 1 0 4784 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_44
timestamp 1666464484
transform 1 0 5152 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_46
timestamp 1666464484
transform 1 0 5336 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_58
timestamp 1666464484
transform 1 0 6440 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_70
timestamp 1666464484
transform 1 0 7544 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_74
timestamp 1666464484
transform 1 0 7912 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_76
timestamp 1666464484
transform 1 0 8096 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_88
timestamp 1666464484
transform 1 0 9200 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_100
timestamp 1666464484
transform 1 0 10304 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_104
timestamp 1666464484
transform 1 0 10672 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_106
timestamp 1666464484
transform 1 0 10856 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_118
timestamp 1666464484
transform 1 0 11960 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_130
timestamp 1666464484
transform 1 0 13064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_134
timestamp 1666464484
transform 1 0 13432 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_136
timestamp 1666464484
transform 1 0 13616 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_148
timestamp 1666464484
transform 1 0 14720 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_160
timestamp 1666464484
transform 1 0 15824 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_164
timestamp 1666464484
transform 1 0 16192 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_166
timestamp 1666464484
transform 1 0 16376 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_178
timestamp 1666464484
transform 1 0 17480 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_190
timestamp 1666464484
transform 1 0 18584 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_194
timestamp 1666464484
transform 1 0 18952 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_196
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_208
timestamp 1666464484
transform 1 0 20240 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_220
timestamp 1666464484
transform 1 0 21344 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_224
timestamp 1666464484
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_226
timestamp 1666464484
transform 1 0 21896 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_238
timestamp 1666464484
transform 1 0 23000 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_250
timestamp 1666464484
transform 1 0 24104 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_254
timestamp 1666464484
transform 1 0 24472 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_256
timestamp 1666464484
transform 1 0 24656 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_268
timestamp 1666464484
transform 1 0 25760 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_280
timestamp 1666464484
transform 1 0 26864 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_284
timestamp 1666464484
transform 1 0 27232 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_286
timestamp 1666464484
transform 1 0 27416 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_298
timestamp 1666464484
transform 1 0 28520 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_310
timestamp 1666464484
transform 1 0 29624 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_314
timestamp 1666464484
transform 1 0 29992 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_316
timestamp 1666464484
transform 1 0 30176 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_328
timestamp 1666464484
transform 1 0 31280 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_340
timestamp 1666464484
transform 1 0 32384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_344
timestamp 1666464484
transform 1 0 32752 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_346
timestamp 1666464484
transform 1 0 32936 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_358
timestamp 1666464484
transform 1 0 34040 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_370
timestamp 1666464484
transform 1 0 35144 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_374
timestamp 1666464484
transform 1 0 35512 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_376
timestamp 1666464484
transform 1 0 35696 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_388
timestamp 1666464484
transform 1 0 36800 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_400
timestamp 1666464484
transform 1 0 37904 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_404
timestamp 1666464484
transform 1 0 38272 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_406
timestamp 1666464484
transform 1 0 38456 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_418
timestamp 1666464484
transform 1 0 39560 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_430
timestamp 1666464484
transform 1 0 40664 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_434
timestamp 1666464484
transform 1 0 41032 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_436
timestamp 1666464484
transform 1 0 41216 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_448
timestamp 1666464484
transform 1 0 42320 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_460
timestamp 1666464484
transform 1 0 43424 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_464
timestamp 1666464484
transform 1 0 43792 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_466
timestamp 1666464484
transform 1 0 43976 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_478
timestamp 1666464484
transform 1 0 45080 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_490
timestamp 1666464484
transform 1 0 46184 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_494
timestamp 1666464484
transform 1 0 46552 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_496
timestamp 1666464484
transform 1 0 46736 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_508
timestamp 1666464484
transform 1 0 47840 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_520
timestamp 1666464484
transform 1 0 48944 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_524
timestamp 1666464484
transform 1 0 49312 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_526
timestamp 1666464484
transform 1 0 49496 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_538
timestamp 1666464484
transform 1 0 50600 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_550
timestamp 1666464484
transform 1 0 51704 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_554
timestamp 1666464484
transform 1 0 52072 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_556
timestamp 1666464484
transform 1 0 52256 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_568
timestamp 1666464484
transform 1 0 53360 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_580
timestamp 1666464484
transform 1 0 54464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_584
timestamp 1666464484
transform 1 0 54832 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_586
timestamp 1666464484
transform 1 0 55016 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_598
timestamp 1666464484
transform 1 0 56120 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_610
timestamp 1666464484
transform 1 0 57224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_614
timestamp 1666464484
transform 1 0 57592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_616
timestamp 1666464484
transform 1 0 57776 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_624
timestamp 1666464484
transform 1 0 58512 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_31
timestamp 1666464484
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_43
timestamp 1666464484
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_59
timestamp 1666464484
transform 1 0 6532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_61
timestamp 1666464484
transform 1 0 6716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_73
timestamp 1666464484
transform 1 0 7820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_85
timestamp 1666464484
transform 1 0 8924 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_89
timestamp 1666464484
transform 1 0 9292 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_91
timestamp 1666464484
transform 1 0 9476 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_103
timestamp 1666464484
transform 1 0 10580 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_115
timestamp 1666464484
transform 1 0 11684 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_119
timestamp 1666464484
transform 1 0 12052 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_121
timestamp 1666464484
transform 1 0 12236 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_133
timestamp 1666464484
transform 1 0 13340 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_145
timestamp 1666464484
transform 1 0 14444 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_149
timestamp 1666464484
transform 1 0 14812 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_151
timestamp 1666464484
transform 1 0 14996 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_163
timestamp 1666464484
transform 1 0 16100 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_175
timestamp 1666464484
transform 1 0 17204 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_179
timestamp 1666464484
transform 1 0 17572 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1666464484
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_205
timestamp 1666464484
transform 1 0 19964 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_209
timestamp 1666464484
transform 1 0 20332 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_211
timestamp 1666464484
transform 1 0 20516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_223
timestamp 1666464484
transform 1 0 21620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_235
timestamp 1666464484
transform 1 0 22724 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_239
timestamp 1666464484
transform 1 0 23092 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_241
timestamp 1666464484
transform 1 0 23276 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_253
timestamp 1666464484
transform 1 0 24380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_265
timestamp 1666464484
transform 1 0 25484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_269
timestamp 1666464484
transform 1 0 25852 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_271
timestamp 1666464484
transform 1 0 26036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_283
timestamp 1666464484
transform 1 0 27140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_295
timestamp 1666464484
transform 1 0 28244 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_299
timestamp 1666464484
transform 1 0 28612 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_301
timestamp 1666464484
transform 1 0 28796 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_313
timestamp 1666464484
transform 1 0 29900 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_325
timestamp 1666464484
transform 1 0 31004 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_329
timestamp 1666464484
transform 1 0 31372 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_331
timestamp 1666464484
transform 1 0 31556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_343
timestamp 1666464484
transform 1 0 32660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_355
timestamp 1666464484
transform 1 0 33764 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_359
timestamp 1666464484
transform 1 0 34132 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1666464484
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1666464484
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_385
timestamp 1666464484
transform 1 0 36524 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_389
timestamp 1666464484
transform 1 0 36892 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_391
timestamp 1666464484
transform 1 0 37076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_403
timestamp 1666464484
transform 1 0 38180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_415
timestamp 1666464484
transform 1 0 39284 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_419
timestamp 1666464484
transform 1 0 39652 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_421
timestamp 1666464484
transform 1 0 39836 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_433
timestamp 1666464484
transform 1 0 40940 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_445
timestamp 1666464484
transform 1 0 42044 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_449
timestamp 1666464484
transform 1 0 42412 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_451
timestamp 1666464484
transform 1 0 42596 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_463
timestamp 1666464484
transform 1 0 43700 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_475
timestamp 1666464484
transform 1 0 44804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_479
timestamp 1666464484
transform 1 0 45172 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_481
timestamp 1666464484
transform 1 0 45356 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_493
timestamp 1666464484
transform 1 0 46460 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_505
timestamp 1666464484
transform 1 0 47564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_509
timestamp 1666464484
transform 1 0 47932 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_511
timestamp 1666464484
transform 1 0 48116 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_523
timestamp 1666464484
transform 1 0 49220 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_535
timestamp 1666464484
transform 1 0 50324 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_539
timestamp 1666464484
transform 1 0 50692 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1666464484
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_553
timestamp 1666464484
transform 1 0 51980 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_565
timestamp 1666464484
transform 1 0 53084 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_569
timestamp 1666464484
transform 1 0 53452 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_571
timestamp 1666464484
transform 1 0 53636 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_583
timestamp 1666464484
transform 1 0 54740 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_595
timestamp 1666464484
transform 1 0 55844 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_599
timestamp 1666464484
transform 1 0 56212 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_601
timestamp 1666464484
transform 1 0 56396 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_613
timestamp 1666464484
transform 1 0 57500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_16
timestamp 1666464484
transform 1 0 2576 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_28
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_40
timestamp 1666464484
transform 1 0 4784 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_44
timestamp 1666464484
transform 1 0 5152 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_46
timestamp 1666464484
transform 1 0 5336 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_58
timestamp 1666464484
transform 1 0 6440 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_70
timestamp 1666464484
transform 1 0 7544 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_74
timestamp 1666464484
transform 1 0 7912 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_76
timestamp 1666464484
transform 1 0 8096 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_88
timestamp 1666464484
transform 1 0 9200 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_100
timestamp 1666464484
transform 1 0 10304 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_104
timestamp 1666464484
transform 1 0 10672 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_106
timestamp 1666464484
transform 1 0 10856 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_118
timestamp 1666464484
transform 1 0 11960 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_130
timestamp 1666464484
transform 1 0 13064 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_134
timestamp 1666464484
transform 1 0 13432 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_136
timestamp 1666464484
transform 1 0 13616 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_148
timestamp 1666464484
transform 1 0 14720 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_160
timestamp 1666464484
transform 1 0 15824 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_164
timestamp 1666464484
transform 1 0 16192 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_166
timestamp 1666464484
transform 1 0 16376 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_178
timestamp 1666464484
transform 1 0 17480 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_190
timestamp 1666464484
transform 1 0 18584 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_194
timestamp 1666464484
transform 1 0 18952 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_196
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_208
timestamp 1666464484
transform 1 0 20240 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_220
timestamp 1666464484
transform 1 0 21344 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_224
timestamp 1666464484
transform 1 0 21712 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_226
timestamp 1666464484
transform 1 0 21896 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_238
timestamp 1666464484
transform 1 0 23000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_250
timestamp 1666464484
transform 1 0 24104 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_254
timestamp 1666464484
transform 1 0 24472 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_256
timestamp 1666464484
transform 1 0 24656 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_268
timestamp 1666464484
transform 1 0 25760 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_280
timestamp 1666464484
transform 1 0 26864 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_284
timestamp 1666464484
transform 1 0 27232 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_286
timestamp 1666464484
transform 1 0 27416 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_298
timestamp 1666464484
transform 1 0 28520 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_310
timestamp 1666464484
transform 1 0 29624 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_314
timestamp 1666464484
transform 1 0 29992 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_316
timestamp 1666464484
transform 1 0 30176 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_328
timestamp 1666464484
transform 1 0 31280 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_340
timestamp 1666464484
transform 1 0 32384 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_344
timestamp 1666464484
transform 1 0 32752 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_346
timestamp 1666464484
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_358
timestamp 1666464484
transform 1 0 34040 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_370
timestamp 1666464484
transform 1 0 35144 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_374
timestamp 1666464484
transform 1 0 35512 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_376
timestamp 1666464484
transform 1 0 35696 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_388
timestamp 1666464484
transform 1 0 36800 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_400
timestamp 1666464484
transform 1 0 37904 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_404
timestamp 1666464484
transform 1 0 38272 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_406
timestamp 1666464484
transform 1 0 38456 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_418
timestamp 1666464484
transform 1 0 39560 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_430
timestamp 1666464484
transform 1 0 40664 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_434
timestamp 1666464484
transform 1 0 41032 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_436
timestamp 1666464484
transform 1 0 41216 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_448
timestamp 1666464484
transform 1 0 42320 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_460
timestamp 1666464484
transform 1 0 43424 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_464
timestamp 1666464484
transform 1 0 43792 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_466
timestamp 1666464484
transform 1 0 43976 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_478
timestamp 1666464484
transform 1 0 45080 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_490
timestamp 1666464484
transform 1 0 46184 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_494
timestamp 1666464484
transform 1 0 46552 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_496
timestamp 1666464484
transform 1 0 46736 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_508
timestamp 1666464484
transform 1 0 47840 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_520
timestamp 1666464484
transform 1 0 48944 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_524
timestamp 1666464484
transform 1 0 49312 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_526
timestamp 1666464484
transform 1 0 49496 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_538
timestamp 1666464484
transform 1 0 50600 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_550
timestamp 1666464484
transform 1 0 51704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_554
timestamp 1666464484
transform 1 0 52072 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_556
timestamp 1666464484
transform 1 0 52256 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_568
timestamp 1666464484
transform 1 0 53360 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_580
timestamp 1666464484
transform 1 0 54464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_584
timestamp 1666464484
transform 1 0 54832 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_586
timestamp 1666464484
transform 1 0 55016 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_598
timestamp 1666464484
transform 1 0 56120 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_610
timestamp 1666464484
transform 1 0 57224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_614
timestamp 1666464484
transform 1 0 57592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_616
timestamp 1666464484
transform 1 0 57776 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_624
timestamp 1666464484
transform 1 0 58512 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666464484
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_27
timestamp 1666464484
transform 1 0 3588 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_31
timestamp 1666464484
transform 1 0 3956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_43
timestamp 1666464484
transform 1 0 5060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_55
timestamp 1666464484
transform 1 0 6164 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_59
timestamp 1666464484
transform 1 0 6532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_61
timestamp 1666464484
transform 1 0 6716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_73
timestamp 1666464484
transform 1 0 7820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_85
timestamp 1666464484
transform 1 0 8924 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_89
timestamp 1666464484
transform 1 0 9292 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_91
timestamp 1666464484
transform 1 0 9476 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_103
timestamp 1666464484
transform 1 0 10580 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_115
timestamp 1666464484
transform 1 0 11684 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_119
timestamp 1666464484
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_121
timestamp 1666464484
transform 1 0 12236 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_133
timestamp 1666464484
transform 1 0 13340 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_145
timestamp 1666464484
transform 1 0 14444 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_149
timestamp 1666464484
transform 1 0 14812 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_151
timestamp 1666464484
transform 1 0 14996 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_163
timestamp 1666464484
transform 1 0 16100 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_175
timestamp 1666464484
transform 1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_179
timestamp 1666464484
transform 1 0 17572 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1666464484
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_205
timestamp 1666464484
transform 1 0 19964 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_209
timestamp 1666464484
transform 1 0 20332 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_211
timestamp 1666464484
transform 1 0 20516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_223
timestamp 1666464484
transform 1 0 21620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_235
timestamp 1666464484
transform 1 0 22724 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_239
timestamp 1666464484
transform 1 0 23092 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_241
timestamp 1666464484
transform 1 0 23276 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_253
timestamp 1666464484
transform 1 0 24380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_265
timestamp 1666464484
transform 1 0 25484 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_269
timestamp 1666464484
transform 1 0 25852 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_271
timestamp 1666464484
transform 1 0 26036 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_283
timestamp 1666464484
transform 1 0 27140 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_295
timestamp 1666464484
transform 1 0 28244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_299
timestamp 1666464484
transform 1 0 28612 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_301
timestamp 1666464484
transform 1 0 28796 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_313
timestamp 1666464484
transform 1 0 29900 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_325
timestamp 1666464484
transform 1 0 31004 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_329
timestamp 1666464484
transform 1 0 31372 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_331
timestamp 1666464484
transform 1 0 31556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_343
timestamp 1666464484
transform 1 0 32660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_355
timestamp 1666464484
transform 1 0 33764 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_359
timestamp 1666464484
transform 1 0 34132 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1666464484
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1666464484
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_385
timestamp 1666464484
transform 1 0 36524 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_389
timestamp 1666464484
transform 1 0 36892 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_391
timestamp 1666464484
transform 1 0 37076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_403
timestamp 1666464484
transform 1 0 38180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_415
timestamp 1666464484
transform 1 0 39284 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_419
timestamp 1666464484
transform 1 0 39652 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_421
timestamp 1666464484
transform 1 0 39836 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_433
timestamp 1666464484
transform 1 0 40940 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_445
timestamp 1666464484
transform 1 0 42044 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_449
timestamp 1666464484
transform 1 0 42412 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_451
timestamp 1666464484
transform 1 0 42596 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_463
timestamp 1666464484
transform 1 0 43700 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_475
timestamp 1666464484
transform 1 0 44804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_479
timestamp 1666464484
transform 1 0 45172 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_481
timestamp 1666464484
transform 1 0 45356 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_493
timestamp 1666464484
transform 1 0 46460 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_505
timestamp 1666464484
transform 1 0 47564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_509
timestamp 1666464484
transform 1 0 47932 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_511
timestamp 1666464484
transform 1 0 48116 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_523
timestamp 1666464484
transform 1 0 49220 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_535
timestamp 1666464484
transform 1 0 50324 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_539
timestamp 1666464484
transform 1 0 50692 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1666464484
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_553
timestamp 1666464484
transform 1 0 51980 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_565
timestamp 1666464484
transform 1 0 53084 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_569
timestamp 1666464484
transform 1 0 53452 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_571
timestamp 1666464484
transform 1 0 53636 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_583
timestamp 1666464484
transform 1 0 54740 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_595
timestamp 1666464484
transform 1 0 55844 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_599
timestamp 1666464484
transform 1 0 56212 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_601
timestamp 1666464484
transform 1 0 56396 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_613
timestamp 1666464484
transform 1 0 57500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_16
timestamp 1666464484
transform 1 0 2576 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_28
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_40
timestamp 1666464484
transform 1 0 4784 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_44
timestamp 1666464484
transform 1 0 5152 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_46
timestamp 1666464484
transform 1 0 5336 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_58
timestamp 1666464484
transform 1 0 6440 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_70
timestamp 1666464484
transform 1 0 7544 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_74
timestamp 1666464484
transform 1 0 7912 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_76
timestamp 1666464484
transform 1 0 8096 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_88
timestamp 1666464484
transform 1 0 9200 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_100
timestamp 1666464484
transform 1 0 10304 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_104
timestamp 1666464484
transform 1 0 10672 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_106
timestamp 1666464484
transform 1 0 10856 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_118
timestamp 1666464484
transform 1 0 11960 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_130
timestamp 1666464484
transform 1 0 13064 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_134
timestamp 1666464484
transform 1 0 13432 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_136
timestamp 1666464484
transform 1 0 13616 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_148
timestamp 1666464484
transform 1 0 14720 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_160
timestamp 1666464484
transform 1 0 15824 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_164
timestamp 1666464484
transform 1 0 16192 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_166
timestamp 1666464484
transform 1 0 16376 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_178
timestamp 1666464484
transform 1 0 17480 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_190
timestamp 1666464484
transform 1 0 18584 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_194
timestamp 1666464484
transform 1 0 18952 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_196
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_208
timestamp 1666464484
transform 1 0 20240 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_220
timestamp 1666464484
transform 1 0 21344 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_224
timestamp 1666464484
transform 1 0 21712 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_226
timestamp 1666464484
transform 1 0 21896 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_238
timestamp 1666464484
transform 1 0 23000 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_250
timestamp 1666464484
transform 1 0 24104 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_254
timestamp 1666464484
transform 1 0 24472 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_256
timestamp 1666464484
transform 1 0 24656 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_268
timestamp 1666464484
transform 1 0 25760 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_280
timestamp 1666464484
transform 1 0 26864 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_284
timestamp 1666464484
transform 1 0 27232 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_286
timestamp 1666464484
transform 1 0 27416 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_298
timestamp 1666464484
transform 1 0 28520 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_310
timestamp 1666464484
transform 1 0 29624 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_314
timestamp 1666464484
transform 1 0 29992 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_316
timestamp 1666464484
transform 1 0 30176 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_328
timestamp 1666464484
transform 1 0 31280 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_340
timestamp 1666464484
transform 1 0 32384 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_344
timestamp 1666464484
transform 1 0 32752 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_346
timestamp 1666464484
transform 1 0 32936 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_358
timestamp 1666464484
transform 1 0 34040 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_370
timestamp 1666464484
transform 1 0 35144 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_374
timestamp 1666464484
transform 1 0 35512 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_376
timestamp 1666464484
transform 1 0 35696 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_388
timestamp 1666464484
transform 1 0 36800 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_400
timestamp 1666464484
transform 1 0 37904 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_404
timestamp 1666464484
transform 1 0 38272 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_406
timestamp 1666464484
transform 1 0 38456 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_418
timestamp 1666464484
transform 1 0 39560 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_430
timestamp 1666464484
transform 1 0 40664 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_434
timestamp 1666464484
transform 1 0 41032 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_436
timestamp 1666464484
transform 1 0 41216 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_448
timestamp 1666464484
transform 1 0 42320 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_460
timestamp 1666464484
transform 1 0 43424 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_464
timestamp 1666464484
transform 1 0 43792 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_466
timestamp 1666464484
transform 1 0 43976 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_478
timestamp 1666464484
transform 1 0 45080 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_490
timestamp 1666464484
transform 1 0 46184 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_494
timestamp 1666464484
transform 1 0 46552 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_496
timestamp 1666464484
transform 1 0 46736 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_508
timestamp 1666464484
transform 1 0 47840 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_520
timestamp 1666464484
transform 1 0 48944 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_524
timestamp 1666464484
transform 1 0 49312 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_526
timestamp 1666464484
transform 1 0 49496 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_538
timestamp 1666464484
transform 1 0 50600 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_550
timestamp 1666464484
transform 1 0 51704 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_554
timestamp 1666464484
transform 1 0 52072 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_556
timestamp 1666464484
transform 1 0 52256 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_568
timestamp 1666464484
transform 1 0 53360 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_580
timestamp 1666464484
transform 1 0 54464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_584
timestamp 1666464484
transform 1 0 54832 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_586
timestamp 1666464484
transform 1 0 55016 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_598
timestamp 1666464484
transform 1 0 56120 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_610
timestamp 1666464484
transform 1 0 57224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_614
timestamp 1666464484
transform 1 0 57592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_616
timestamp 1666464484
transform 1 0 57776 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_624
timestamp 1666464484
transform 1 0 58512 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_31
timestamp 1666464484
transform 1 0 3956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_43
timestamp 1666464484
transform 1 0 5060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_59
timestamp 1666464484
transform 1 0 6532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_61
timestamp 1666464484
transform 1 0 6716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_73
timestamp 1666464484
transform 1 0 7820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_85
timestamp 1666464484
transform 1 0 8924 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_89
timestamp 1666464484
transform 1 0 9292 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_91
timestamp 1666464484
transform 1 0 9476 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_103
timestamp 1666464484
transform 1 0 10580 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_115
timestamp 1666464484
transform 1 0 11684 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_119
timestamp 1666464484
transform 1 0 12052 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_121
timestamp 1666464484
transform 1 0 12236 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_133
timestamp 1666464484
transform 1 0 13340 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_145
timestamp 1666464484
transform 1 0 14444 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_149
timestamp 1666464484
transform 1 0 14812 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_151
timestamp 1666464484
transform 1 0 14996 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_163
timestamp 1666464484
transform 1 0 16100 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_175
timestamp 1666464484
transform 1 0 17204 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_179
timestamp 1666464484
transform 1 0 17572 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1666464484
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1666464484
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_205
timestamp 1666464484
transform 1 0 19964 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_209
timestamp 1666464484
transform 1 0 20332 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_211
timestamp 1666464484
transform 1 0 20516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_223
timestamp 1666464484
transform 1 0 21620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_235
timestamp 1666464484
transform 1 0 22724 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_239
timestamp 1666464484
transform 1 0 23092 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_241
timestamp 1666464484
transform 1 0 23276 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_253
timestamp 1666464484
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_265
timestamp 1666464484
transform 1 0 25484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_269
timestamp 1666464484
transform 1 0 25852 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_271
timestamp 1666464484
transform 1 0 26036 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_283
timestamp 1666464484
transform 1 0 27140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_295
timestamp 1666464484
transform 1 0 28244 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_299
timestamp 1666464484
transform 1 0 28612 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_301
timestamp 1666464484
transform 1 0 28796 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_313
timestamp 1666464484
transform 1 0 29900 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_325
timestamp 1666464484
transform 1 0 31004 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_329
timestamp 1666464484
transform 1 0 31372 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_331
timestamp 1666464484
transform 1 0 31556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_343
timestamp 1666464484
transform 1 0 32660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_355
timestamp 1666464484
transform 1 0 33764 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_359
timestamp 1666464484
transform 1 0 34132 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1666464484
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1666464484
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_385
timestamp 1666464484
transform 1 0 36524 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_389
timestamp 1666464484
transform 1 0 36892 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_391
timestamp 1666464484
transform 1 0 37076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_403
timestamp 1666464484
transform 1 0 38180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_415
timestamp 1666464484
transform 1 0 39284 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_419
timestamp 1666464484
transform 1 0 39652 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_421
timestamp 1666464484
transform 1 0 39836 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_433
timestamp 1666464484
transform 1 0 40940 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_445
timestamp 1666464484
transform 1 0 42044 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_449
timestamp 1666464484
transform 1 0 42412 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_451
timestamp 1666464484
transform 1 0 42596 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_463
timestamp 1666464484
transform 1 0 43700 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_475
timestamp 1666464484
transform 1 0 44804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_479
timestamp 1666464484
transform 1 0 45172 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_481
timestamp 1666464484
transform 1 0 45356 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_493
timestamp 1666464484
transform 1 0 46460 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_505
timestamp 1666464484
transform 1 0 47564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_509
timestamp 1666464484
transform 1 0 47932 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_511
timestamp 1666464484
transform 1 0 48116 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_523
timestamp 1666464484
transform 1 0 49220 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_535
timestamp 1666464484
transform 1 0 50324 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_539
timestamp 1666464484
transform 1 0 50692 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1666464484
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_553
timestamp 1666464484
transform 1 0 51980 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_565
timestamp 1666464484
transform 1 0 53084 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_569
timestamp 1666464484
transform 1 0 53452 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_571
timestamp 1666464484
transform 1 0 53636 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_583
timestamp 1666464484
transform 1 0 54740 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_595
timestamp 1666464484
transform 1 0 55844 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_599
timestamp 1666464484
transform 1 0 56212 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_601
timestamp 1666464484
transform 1 0 56396 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_613
timestamp 1666464484
transform 1 0 57500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_16
timestamp 1666464484
transform 1 0 2576 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_28
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_40
timestamp 1666464484
transform 1 0 4784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_44
timestamp 1666464484
transform 1 0 5152 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_46
timestamp 1666464484
transform 1 0 5336 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_58
timestamp 1666464484
transform 1 0 6440 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_70
timestamp 1666464484
transform 1 0 7544 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_74
timestamp 1666464484
transform 1 0 7912 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_76
timestamp 1666464484
transform 1 0 8096 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_88
timestamp 1666464484
transform 1 0 9200 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_100
timestamp 1666464484
transform 1 0 10304 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_104
timestamp 1666464484
transform 1 0 10672 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_106
timestamp 1666464484
transform 1 0 10856 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_118
timestamp 1666464484
transform 1 0 11960 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_130
timestamp 1666464484
transform 1 0 13064 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_134
timestamp 1666464484
transform 1 0 13432 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_136
timestamp 1666464484
transform 1 0 13616 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_148
timestamp 1666464484
transform 1 0 14720 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_160
timestamp 1666464484
transform 1 0 15824 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_164
timestamp 1666464484
transform 1 0 16192 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_166
timestamp 1666464484
transform 1 0 16376 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_178
timestamp 1666464484
transform 1 0 17480 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_190
timestamp 1666464484
transform 1 0 18584 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_194
timestamp 1666464484
transform 1 0 18952 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_196
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_208
timestamp 1666464484
transform 1 0 20240 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_220
timestamp 1666464484
transform 1 0 21344 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_224
timestamp 1666464484
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_226
timestamp 1666464484
transform 1 0 21896 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_238
timestamp 1666464484
transform 1 0 23000 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_250
timestamp 1666464484
transform 1 0 24104 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_254
timestamp 1666464484
transform 1 0 24472 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_256
timestamp 1666464484
transform 1 0 24656 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_268
timestamp 1666464484
transform 1 0 25760 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_280
timestamp 1666464484
transform 1 0 26864 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_284
timestamp 1666464484
transform 1 0 27232 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_286
timestamp 1666464484
transform 1 0 27416 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_298
timestamp 1666464484
transform 1 0 28520 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_310
timestamp 1666464484
transform 1 0 29624 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_314
timestamp 1666464484
transform 1 0 29992 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_316
timestamp 1666464484
transform 1 0 30176 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_328
timestamp 1666464484
transform 1 0 31280 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_340
timestamp 1666464484
transform 1 0 32384 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_344
timestamp 1666464484
transform 1 0 32752 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_346
timestamp 1666464484
transform 1 0 32936 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_358
timestamp 1666464484
transform 1 0 34040 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_370
timestamp 1666464484
transform 1 0 35144 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_374
timestamp 1666464484
transform 1 0 35512 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_376
timestamp 1666464484
transform 1 0 35696 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_388
timestamp 1666464484
transform 1 0 36800 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_400
timestamp 1666464484
transform 1 0 37904 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_404
timestamp 1666464484
transform 1 0 38272 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_406
timestamp 1666464484
transform 1 0 38456 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_418
timestamp 1666464484
transform 1 0 39560 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_430
timestamp 1666464484
transform 1 0 40664 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_434
timestamp 1666464484
transform 1 0 41032 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_436
timestamp 1666464484
transform 1 0 41216 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_448
timestamp 1666464484
transform 1 0 42320 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_460
timestamp 1666464484
transform 1 0 43424 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_464
timestamp 1666464484
transform 1 0 43792 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_466
timestamp 1666464484
transform 1 0 43976 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_478
timestamp 1666464484
transform 1 0 45080 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_490
timestamp 1666464484
transform 1 0 46184 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_494
timestamp 1666464484
transform 1 0 46552 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_496
timestamp 1666464484
transform 1 0 46736 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_508
timestamp 1666464484
transform 1 0 47840 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_520
timestamp 1666464484
transform 1 0 48944 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_524
timestamp 1666464484
transform 1 0 49312 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_526
timestamp 1666464484
transform 1 0 49496 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_538
timestamp 1666464484
transform 1 0 50600 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_550
timestamp 1666464484
transform 1 0 51704 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_554
timestamp 1666464484
transform 1 0 52072 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_556
timestamp 1666464484
transform 1 0 52256 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_568
timestamp 1666464484
transform 1 0 53360 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_580
timestamp 1666464484
transform 1 0 54464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_584
timestamp 1666464484
transform 1 0 54832 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_586
timestamp 1666464484
transform 1 0 55016 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_598
timestamp 1666464484
transform 1 0 56120 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_610
timestamp 1666464484
transform 1 0 57224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_614
timestamp 1666464484
transform 1 0 57592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_616
timestamp 1666464484
transform 1 0 57776 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_624
timestamp 1666464484
transform 1 0 58512 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_31
timestamp 1666464484
transform 1 0 3956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_43
timestamp 1666464484
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_55
timestamp 1666464484
transform 1 0 6164 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_59
timestamp 1666464484
transform 1 0 6532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_61
timestamp 1666464484
transform 1 0 6716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_73
timestamp 1666464484
transform 1 0 7820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_85
timestamp 1666464484
transform 1 0 8924 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_89
timestamp 1666464484
transform 1 0 9292 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_91
timestamp 1666464484
transform 1 0 9476 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_103
timestamp 1666464484
transform 1 0 10580 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_115
timestamp 1666464484
transform 1 0 11684 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_119
timestamp 1666464484
transform 1 0 12052 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_121
timestamp 1666464484
transform 1 0 12236 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_133
timestamp 1666464484
transform 1 0 13340 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_145
timestamp 1666464484
transform 1 0 14444 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_149
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_151
timestamp 1666464484
transform 1 0 14996 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_163
timestamp 1666464484
transform 1 0 16100 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_175
timestamp 1666464484
transform 1 0 17204 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_179
timestamp 1666464484
transform 1 0 17572 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666464484
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1666464484
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_205
timestamp 1666464484
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_209
timestamp 1666464484
transform 1 0 20332 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_211
timestamp 1666464484
transform 1 0 20516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_223
timestamp 1666464484
transform 1 0 21620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_235
timestamp 1666464484
transform 1 0 22724 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_239
timestamp 1666464484
transform 1 0 23092 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_241
timestamp 1666464484
transform 1 0 23276 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_253
timestamp 1666464484
transform 1 0 24380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_265
timestamp 1666464484
transform 1 0 25484 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_269
timestamp 1666464484
transform 1 0 25852 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_271
timestamp 1666464484
transform 1 0 26036 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_283
timestamp 1666464484
transform 1 0 27140 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_295
timestamp 1666464484
transform 1 0 28244 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_299
timestamp 1666464484
transform 1 0 28612 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_301
timestamp 1666464484
transform 1 0 28796 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_313
timestamp 1666464484
transform 1 0 29900 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_325
timestamp 1666464484
transform 1 0 31004 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_329
timestamp 1666464484
transform 1 0 31372 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_331
timestamp 1666464484
transform 1 0 31556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_343
timestamp 1666464484
transform 1 0 32660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_355
timestamp 1666464484
transform 1 0 33764 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_359
timestamp 1666464484
transform 1 0 34132 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1666464484
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1666464484
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_385
timestamp 1666464484
transform 1 0 36524 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_389
timestamp 1666464484
transform 1 0 36892 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_391
timestamp 1666464484
transform 1 0 37076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_403
timestamp 1666464484
transform 1 0 38180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_415
timestamp 1666464484
transform 1 0 39284 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_419
timestamp 1666464484
transform 1 0 39652 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_421
timestamp 1666464484
transform 1 0 39836 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_433
timestamp 1666464484
transform 1 0 40940 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_445
timestamp 1666464484
transform 1 0 42044 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_449
timestamp 1666464484
transform 1 0 42412 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_451
timestamp 1666464484
transform 1 0 42596 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_463
timestamp 1666464484
transform 1 0 43700 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_475
timestamp 1666464484
transform 1 0 44804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_479
timestamp 1666464484
transform 1 0 45172 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_481
timestamp 1666464484
transform 1 0 45356 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_493
timestamp 1666464484
transform 1 0 46460 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_505
timestamp 1666464484
transform 1 0 47564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_509
timestamp 1666464484
transform 1 0 47932 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_511
timestamp 1666464484
transform 1 0 48116 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_523
timestamp 1666464484
transform 1 0 49220 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_535
timestamp 1666464484
transform 1 0 50324 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_539
timestamp 1666464484
transform 1 0 50692 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1666464484
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_553
timestamp 1666464484
transform 1 0 51980 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_565
timestamp 1666464484
transform 1 0 53084 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_569
timestamp 1666464484
transform 1 0 53452 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_571
timestamp 1666464484
transform 1 0 53636 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_583
timestamp 1666464484
transform 1 0 54740 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_595
timestamp 1666464484
transform 1 0 55844 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_599
timestamp 1666464484
transform 1 0 56212 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_601
timestamp 1666464484
transform 1 0 56396 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_613
timestamp 1666464484
transform 1 0 57500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_16
timestamp 1666464484
transform 1 0 2576 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_28
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_40
timestamp 1666464484
transform 1 0 4784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_44
timestamp 1666464484
transform 1 0 5152 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_46
timestamp 1666464484
transform 1 0 5336 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_58
timestamp 1666464484
transform 1 0 6440 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_70
timestamp 1666464484
transform 1 0 7544 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_74
timestamp 1666464484
transform 1 0 7912 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_76
timestamp 1666464484
transform 1 0 8096 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_88
timestamp 1666464484
transform 1 0 9200 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_100
timestamp 1666464484
transform 1 0 10304 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_104
timestamp 1666464484
transform 1 0 10672 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_106
timestamp 1666464484
transform 1 0 10856 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_118
timestamp 1666464484
transform 1 0 11960 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_130
timestamp 1666464484
transform 1 0 13064 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_134
timestamp 1666464484
transform 1 0 13432 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_136
timestamp 1666464484
transform 1 0 13616 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_148
timestamp 1666464484
transform 1 0 14720 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_160
timestamp 1666464484
transform 1 0 15824 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_164
timestamp 1666464484
transform 1 0 16192 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_166
timestamp 1666464484
transform 1 0 16376 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_178
timestamp 1666464484
transform 1 0 17480 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_190
timestamp 1666464484
transform 1 0 18584 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_194
timestamp 1666464484
transform 1 0 18952 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_196
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_208
timestamp 1666464484
transform 1 0 20240 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_220
timestamp 1666464484
transform 1 0 21344 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_224
timestamp 1666464484
transform 1 0 21712 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_226
timestamp 1666464484
transform 1 0 21896 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_238
timestamp 1666464484
transform 1 0 23000 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_250
timestamp 1666464484
transform 1 0 24104 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_254
timestamp 1666464484
transform 1 0 24472 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_256
timestamp 1666464484
transform 1 0 24656 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_268
timestamp 1666464484
transform 1 0 25760 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_280
timestamp 1666464484
transform 1 0 26864 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_284
timestamp 1666464484
transform 1 0 27232 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_286
timestamp 1666464484
transform 1 0 27416 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_298
timestamp 1666464484
transform 1 0 28520 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_310
timestamp 1666464484
transform 1 0 29624 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_314
timestamp 1666464484
transform 1 0 29992 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_316
timestamp 1666464484
transform 1 0 30176 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_328
timestamp 1666464484
transform 1 0 31280 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_340
timestamp 1666464484
transform 1 0 32384 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_344
timestamp 1666464484
transform 1 0 32752 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_346
timestamp 1666464484
transform 1 0 32936 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_358
timestamp 1666464484
transform 1 0 34040 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_370
timestamp 1666464484
transform 1 0 35144 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_374
timestamp 1666464484
transform 1 0 35512 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_376
timestamp 1666464484
transform 1 0 35696 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_388
timestamp 1666464484
transform 1 0 36800 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_400
timestamp 1666464484
transform 1 0 37904 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_404
timestamp 1666464484
transform 1 0 38272 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_406
timestamp 1666464484
transform 1 0 38456 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_418
timestamp 1666464484
transform 1 0 39560 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_430
timestamp 1666464484
transform 1 0 40664 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_434
timestamp 1666464484
transform 1 0 41032 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_436
timestamp 1666464484
transform 1 0 41216 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_448
timestamp 1666464484
transform 1 0 42320 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_460
timestamp 1666464484
transform 1 0 43424 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_464
timestamp 1666464484
transform 1 0 43792 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_466
timestamp 1666464484
transform 1 0 43976 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_478
timestamp 1666464484
transform 1 0 45080 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_490
timestamp 1666464484
transform 1 0 46184 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_494
timestamp 1666464484
transform 1 0 46552 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_496
timestamp 1666464484
transform 1 0 46736 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_508
timestamp 1666464484
transform 1 0 47840 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_520
timestamp 1666464484
transform 1 0 48944 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_524
timestamp 1666464484
transform 1 0 49312 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_526
timestamp 1666464484
transform 1 0 49496 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_538
timestamp 1666464484
transform 1 0 50600 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_550
timestamp 1666464484
transform 1 0 51704 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_554
timestamp 1666464484
transform 1 0 52072 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_556
timestamp 1666464484
transform 1 0 52256 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_568
timestamp 1666464484
transform 1 0 53360 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_580
timestamp 1666464484
transform 1 0 54464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_584
timestamp 1666464484
transform 1 0 54832 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_586
timestamp 1666464484
transform 1 0 55016 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_598
timestamp 1666464484
transform 1 0 56120 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_610
timestamp 1666464484
transform 1 0 57224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_614
timestamp 1666464484
transform 1 0 57592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_616
timestamp 1666464484
transform 1 0 57776 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_624
timestamp 1666464484
transform 1 0 58512 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_31
timestamp 1666464484
transform 1 0 3956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_43
timestamp 1666464484
transform 1 0 5060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_59
timestamp 1666464484
transform 1 0 6532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_61
timestamp 1666464484
transform 1 0 6716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_73
timestamp 1666464484
transform 1 0 7820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_85
timestamp 1666464484
transform 1 0 8924 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_89
timestamp 1666464484
transform 1 0 9292 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_91
timestamp 1666464484
transform 1 0 9476 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_103
timestamp 1666464484
transform 1 0 10580 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_115
timestamp 1666464484
transform 1 0 11684 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_119
timestamp 1666464484
transform 1 0 12052 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_121
timestamp 1666464484
transform 1 0 12236 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_133
timestamp 1666464484
transform 1 0 13340 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_145
timestamp 1666464484
transform 1 0 14444 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_149
timestamp 1666464484
transform 1 0 14812 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_151
timestamp 1666464484
transform 1 0 14996 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_163
timestamp 1666464484
transform 1 0 16100 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_175
timestamp 1666464484
transform 1 0 17204 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_179
timestamp 1666464484
transform 1 0 17572 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1666464484
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1666464484
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_205
timestamp 1666464484
transform 1 0 19964 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_209
timestamp 1666464484
transform 1 0 20332 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_211
timestamp 1666464484
transform 1 0 20516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_223
timestamp 1666464484
transform 1 0 21620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_235
timestamp 1666464484
transform 1 0 22724 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_239
timestamp 1666464484
transform 1 0 23092 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_241
timestamp 1666464484
transform 1 0 23276 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_253
timestamp 1666464484
transform 1 0 24380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_265
timestamp 1666464484
transform 1 0 25484 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_269
timestamp 1666464484
transform 1 0 25852 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_271
timestamp 1666464484
transform 1 0 26036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_283
timestamp 1666464484
transform 1 0 27140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_295
timestamp 1666464484
transform 1 0 28244 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_299
timestamp 1666464484
transform 1 0 28612 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_301
timestamp 1666464484
transform 1 0 28796 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_313
timestamp 1666464484
transform 1 0 29900 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_325
timestamp 1666464484
transform 1 0 31004 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_329
timestamp 1666464484
transform 1 0 31372 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_331
timestamp 1666464484
transform 1 0 31556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_343
timestamp 1666464484
transform 1 0 32660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_355
timestamp 1666464484
transform 1 0 33764 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_359
timestamp 1666464484
transform 1 0 34132 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1666464484
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1666464484
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_385
timestamp 1666464484
transform 1 0 36524 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_389
timestamp 1666464484
transform 1 0 36892 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_391
timestamp 1666464484
transform 1 0 37076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_403
timestamp 1666464484
transform 1 0 38180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_415
timestamp 1666464484
transform 1 0 39284 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_419
timestamp 1666464484
transform 1 0 39652 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_421
timestamp 1666464484
transform 1 0 39836 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_433
timestamp 1666464484
transform 1 0 40940 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_445
timestamp 1666464484
transform 1 0 42044 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_449
timestamp 1666464484
transform 1 0 42412 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_451
timestamp 1666464484
transform 1 0 42596 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_463
timestamp 1666464484
transform 1 0 43700 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_475
timestamp 1666464484
transform 1 0 44804 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_479
timestamp 1666464484
transform 1 0 45172 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_481
timestamp 1666464484
transform 1 0 45356 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_493
timestamp 1666464484
transform 1 0 46460 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_505
timestamp 1666464484
transform 1 0 47564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_509
timestamp 1666464484
transform 1 0 47932 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_511
timestamp 1666464484
transform 1 0 48116 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_523
timestamp 1666464484
transform 1 0 49220 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_535
timestamp 1666464484
transform 1 0 50324 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_539
timestamp 1666464484
transform 1 0 50692 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1666464484
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_553
timestamp 1666464484
transform 1 0 51980 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_565
timestamp 1666464484
transform 1 0 53084 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_569
timestamp 1666464484
transform 1 0 53452 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_571
timestamp 1666464484
transform 1 0 53636 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_583
timestamp 1666464484
transform 1 0 54740 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_595
timestamp 1666464484
transform 1 0 55844 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_599
timestamp 1666464484
transform 1 0 56212 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_601
timestamp 1666464484
transform 1 0 56396 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_613
timestamp 1666464484
transform 1 0 57500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_16
timestamp 1666464484
transform 1 0 2576 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_28
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_40
timestamp 1666464484
transform 1 0 4784 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_44
timestamp 1666464484
transform 1 0 5152 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_46
timestamp 1666464484
transform 1 0 5336 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_58
timestamp 1666464484
transform 1 0 6440 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_70
timestamp 1666464484
transform 1 0 7544 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_74
timestamp 1666464484
transform 1 0 7912 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_76
timestamp 1666464484
transform 1 0 8096 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_88
timestamp 1666464484
transform 1 0 9200 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_100
timestamp 1666464484
transform 1 0 10304 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_104
timestamp 1666464484
transform 1 0 10672 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_106
timestamp 1666464484
transform 1 0 10856 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_118
timestamp 1666464484
transform 1 0 11960 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_130
timestamp 1666464484
transform 1 0 13064 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_134
timestamp 1666464484
transform 1 0 13432 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_136
timestamp 1666464484
transform 1 0 13616 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_148
timestamp 1666464484
transform 1 0 14720 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_160
timestamp 1666464484
transform 1 0 15824 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_164
timestamp 1666464484
transform 1 0 16192 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_166
timestamp 1666464484
transform 1 0 16376 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_178
timestamp 1666464484
transform 1 0 17480 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_190
timestamp 1666464484
transform 1 0 18584 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_194
timestamp 1666464484
transform 1 0 18952 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_196
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_208
timestamp 1666464484
transform 1 0 20240 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_220
timestamp 1666464484
transform 1 0 21344 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_224
timestamp 1666464484
transform 1 0 21712 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_226
timestamp 1666464484
transform 1 0 21896 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_238
timestamp 1666464484
transform 1 0 23000 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_250
timestamp 1666464484
transform 1 0 24104 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_254
timestamp 1666464484
transform 1 0 24472 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_256
timestamp 1666464484
transform 1 0 24656 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_268
timestamp 1666464484
transform 1 0 25760 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_280
timestamp 1666464484
transform 1 0 26864 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_284
timestamp 1666464484
transform 1 0 27232 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_286
timestamp 1666464484
transform 1 0 27416 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_298
timestamp 1666464484
transform 1 0 28520 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_310
timestamp 1666464484
transform 1 0 29624 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_314
timestamp 1666464484
transform 1 0 29992 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_316
timestamp 1666464484
transform 1 0 30176 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_328
timestamp 1666464484
transform 1 0 31280 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_340
timestamp 1666464484
transform 1 0 32384 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_344
timestamp 1666464484
transform 1 0 32752 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_346
timestamp 1666464484
transform 1 0 32936 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_358
timestamp 1666464484
transform 1 0 34040 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_370
timestamp 1666464484
transform 1 0 35144 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_374
timestamp 1666464484
transform 1 0 35512 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_376
timestamp 1666464484
transform 1 0 35696 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_388
timestamp 1666464484
transform 1 0 36800 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_400
timestamp 1666464484
transform 1 0 37904 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_404
timestamp 1666464484
transform 1 0 38272 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_406
timestamp 1666464484
transform 1 0 38456 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_418
timestamp 1666464484
transform 1 0 39560 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_430
timestamp 1666464484
transform 1 0 40664 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_434
timestamp 1666464484
transform 1 0 41032 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_436
timestamp 1666464484
transform 1 0 41216 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_448
timestamp 1666464484
transform 1 0 42320 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_460
timestamp 1666464484
transform 1 0 43424 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_464
timestamp 1666464484
transform 1 0 43792 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_466
timestamp 1666464484
transform 1 0 43976 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_478
timestamp 1666464484
transform 1 0 45080 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_490
timestamp 1666464484
transform 1 0 46184 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_494
timestamp 1666464484
transform 1 0 46552 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_496
timestamp 1666464484
transform 1 0 46736 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_508
timestamp 1666464484
transform 1 0 47840 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_520
timestamp 1666464484
transform 1 0 48944 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_524
timestamp 1666464484
transform 1 0 49312 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_526
timestamp 1666464484
transform 1 0 49496 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_538
timestamp 1666464484
transform 1 0 50600 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_550
timestamp 1666464484
transform 1 0 51704 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_554
timestamp 1666464484
transform 1 0 52072 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_556
timestamp 1666464484
transform 1 0 52256 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_568
timestamp 1666464484
transform 1 0 53360 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_580
timestamp 1666464484
transform 1 0 54464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_584
timestamp 1666464484
transform 1 0 54832 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_586
timestamp 1666464484
transform 1 0 55016 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_598
timestamp 1666464484
transform 1 0 56120 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_610
timestamp 1666464484
transform 1 0 57224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_614
timestamp 1666464484
transform 1 0 57592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_616
timestamp 1666464484
transform 1 0 57776 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_624
timestamp 1666464484
transform 1 0 58512 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_31
timestamp 1666464484
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_43
timestamp 1666464484
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_59
timestamp 1666464484
transform 1 0 6532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_61
timestamp 1666464484
transform 1 0 6716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_73
timestamp 1666464484
transform 1 0 7820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_85
timestamp 1666464484
transform 1 0 8924 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_89
timestamp 1666464484
transform 1 0 9292 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_91
timestamp 1666464484
transform 1 0 9476 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_103
timestamp 1666464484
transform 1 0 10580 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_115
timestamp 1666464484
transform 1 0 11684 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_119
timestamp 1666464484
transform 1 0 12052 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_121
timestamp 1666464484
transform 1 0 12236 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_133
timestamp 1666464484
transform 1 0 13340 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_145
timestamp 1666464484
transform 1 0 14444 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_149
timestamp 1666464484
transform 1 0 14812 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_151
timestamp 1666464484
transform 1 0 14996 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_163
timestamp 1666464484
transform 1 0 16100 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_175
timestamp 1666464484
transform 1 0 17204 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_179
timestamp 1666464484
transform 1 0 17572 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1666464484
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1666464484
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_205
timestamp 1666464484
transform 1 0 19964 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_209
timestamp 1666464484
transform 1 0 20332 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_211
timestamp 1666464484
transform 1 0 20516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_223
timestamp 1666464484
transform 1 0 21620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_235
timestamp 1666464484
transform 1 0 22724 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_239
timestamp 1666464484
transform 1 0 23092 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_241
timestamp 1666464484
transform 1 0 23276 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_253
timestamp 1666464484
transform 1 0 24380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_265
timestamp 1666464484
transform 1 0 25484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_269
timestamp 1666464484
transform 1 0 25852 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_271
timestamp 1666464484
transform 1 0 26036 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_283
timestamp 1666464484
transform 1 0 27140 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_295
timestamp 1666464484
transform 1 0 28244 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_299
timestamp 1666464484
transform 1 0 28612 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_301
timestamp 1666464484
transform 1 0 28796 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_313
timestamp 1666464484
transform 1 0 29900 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_325
timestamp 1666464484
transform 1 0 31004 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_329
timestamp 1666464484
transform 1 0 31372 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_331
timestamp 1666464484
transform 1 0 31556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_343
timestamp 1666464484
transform 1 0 32660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_355
timestamp 1666464484
transform 1 0 33764 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_359
timestamp 1666464484
transform 1 0 34132 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1666464484
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1666464484
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_385
timestamp 1666464484
transform 1 0 36524 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_389
timestamp 1666464484
transform 1 0 36892 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_391
timestamp 1666464484
transform 1 0 37076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_403
timestamp 1666464484
transform 1 0 38180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_415
timestamp 1666464484
transform 1 0 39284 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_419
timestamp 1666464484
transform 1 0 39652 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_421
timestamp 1666464484
transform 1 0 39836 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_433
timestamp 1666464484
transform 1 0 40940 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_445
timestamp 1666464484
transform 1 0 42044 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_449
timestamp 1666464484
transform 1 0 42412 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_451
timestamp 1666464484
transform 1 0 42596 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_463
timestamp 1666464484
transform 1 0 43700 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_475
timestamp 1666464484
transform 1 0 44804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_479
timestamp 1666464484
transform 1 0 45172 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_481
timestamp 1666464484
transform 1 0 45356 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_493
timestamp 1666464484
transform 1 0 46460 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_505
timestamp 1666464484
transform 1 0 47564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_509
timestamp 1666464484
transform 1 0 47932 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_511
timestamp 1666464484
transform 1 0 48116 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_523
timestamp 1666464484
transform 1 0 49220 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_535
timestamp 1666464484
transform 1 0 50324 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_539
timestamp 1666464484
transform 1 0 50692 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1666464484
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_553
timestamp 1666464484
transform 1 0 51980 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_565
timestamp 1666464484
transform 1 0 53084 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_569
timestamp 1666464484
transform 1 0 53452 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_571
timestamp 1666464484
transform 1 0 53636 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_583
timestamp 1666464484
transform 1 0 54740 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_595
timestamp 1666464484
transform 1 0 55844 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_599
timestamp 1666464484
transform 1 0 56212 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_601
timestamp 1666464484
transform 1 0 56396 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_613
timestamp 1666464484
transform 1 0 57500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_16
timestamp 1666464484
transform 1 0 2576 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_28
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_40
timestamp 1666464484
transform 1 0 4784 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_44
timestamp 1666464484
transform 1 0 5152 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_46
timestamp 1666464484
transform 1 0 5336 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_58
timestamp 1666464484
transform 1 0 6440 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_70
timestamp 1666464484
transform 1 0 7544 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_74
timestamp 1666464484
transform 1 0 7912 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_76
timestamp 1666464484
transform 1 0 8096 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_88
timestamp 1666464484
transform 1 0 9200 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_100
timestamp 1666464484
transform 1 0 10304 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_104
timestamp 1666464484
transform 1 0 10672 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_106
timestamp 1666464484
transform 1 0 10856 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_118
timestamp 1666464484
transform 1 0 11960 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_130
timestamp 1666464484
transform 1 0 13064 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_134
timestamp 1666464484
transform 1 0 13432 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_136
timestamp 1666464484
transform 1 0 13616 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_148
timestamp 1666464484
transform 1 0 14720 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_160
timestamp 1666464484
transform 1 0 15824 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_164
timestamp 1666464484
transform 1 0 16192 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_166
timestamp 1666464484
transform 1 0 16376 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_178
timestamp 1666464484
transform 1 0 17480 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_190
timestamp 1666464484
transform 1 0 18584 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_194
timestamp 1666464484
transform 1 0 18952 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_196
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_208
timestamp 1666464484
transform 1 0 20240 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_220
timestamp 1666464484
transform 1 0 21344 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_224
timestamp 1666464484
transform 1 0 21712 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_226
timestamp 1666464484
transform 1 0 21896 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_238
timestamp 1666464484
transform 1 0 23000 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_250
timestamp 1666464484
transform 1 0 24104 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_254
timestamp 1666464484
transform 1 0 24472 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_256
timestamp 1666464484
transform 1 0 24656 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_268
timestamp 1666464484
transform 1 0 25760 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_280
timestamp 1666464484
transform 1 0 26864 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_284
timestamp 1666464484
transform 1 0 27232 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_286
timestamp 1666464484
transform 1 0 27416 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_298
timestamp 1666464484
transform 1 0 28520 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_310
timestamp 1666464484
transform 1 0 29624 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_314
timestamp 1666464484
transform 1 0 29992 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_316
timestamp 1666464484
transform 1 0 30176 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_328
timestamp 1666464484
transform 1 0 31280 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_340
timestamp 1666464484
transform 1 0 32384 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_344
timestamp 1666464484
transform 1 0 32752 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_346
timestamp 1666464484
transform 1 0 32936 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_358
timestamp 1666464484
transform 1 0 34040 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_370
timestamp 1666464484
transform 1 0 35144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_374
timestamp 1666464484
transform 1 0 35512 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_376
timestamp 1666464484
transform 1 0 35696 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_388
timestamp 1666464484
transform 1 0 36800 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_400
timestamp 1666464484
transform 1 0 37904 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_404
timestamp 1666464484
transform 1 0 38272 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_406
timestamp 1666464484
transform 1 0 38456 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_418
timestamp 1666464484
transform 1 0 39560 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_430
timestamp 1666464484
transform 1 0 40664 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_434
timestamp 1666464484
transform 1 0 41032 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_436
timestamp 1666464484
transform 1 0 41216 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_448
timestamp 1666464484
transform 1 0 42320 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_460
timestamp 1666464484
transform 1 0 43424 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_464
timestamp 1666464484
transform 1 0 43792 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_466
timestamp 1666464484
transform 1 0 43976 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_478
timestamp 1666464484
transform 1 0 45080 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_490
timestamp 1666464484
transform 1 0 46184 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_494
timestamp 1666464484
transform 1 0 46552 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_496
timestamp 1666464484
transform 1 0 46736 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_508
timestamp 1666464484
transform 1 0 47840 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_520
timestamp 1666464484
transform 1 0 48944 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_524
timestamp 1666464484
transform 1 0 49312 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_526
timestamp 1666464484
transform 1 0 49496 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_538
timestamp 1666464484
transform 1 0 50600 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_550
timestamp 1666464484
transform 1 0 51704 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_554
timestamp 1666464484
transform 1 0 52072 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_556
timestamp 1666464484
transform 1 0 52256 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_568
timestamp 1666464484
transform 1 0 53360 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_580
timestamp 1666464484
transform 1 0 54464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_584
timestamp 1666464484
transform 1 0 54832 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_586
timestamp 1666464484
transform 1 0 55016 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_598
timestamp 1666464484
transform 1 0 56120 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_610
timestamp 1666464484
transform 1 0 57224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_614
timestamp 1666464484
transform 1 0 57592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_616
timestamp 1666464484
transform 1 0 57776 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_624
timestamp 1666464484
transform 1 0 58512 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666464484
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_27
timestamp 1666464484
transform 1 0 3588 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_31
timestamp 1666464484
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_43
timestamp 1666464484
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_55
timestamp 1666464484
transform 1 0 6164 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_59
timestamp 1666464484
transform 1 0 6532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_61
timestamp 1666464484
transform 1 0 6716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_73
timestamp 1666464484
transform 1 0 7820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_85
timestamp 1666464484
transform 1 0 8924 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_89
timestamp 1666464484
transform 1 0 9292 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_91
timestamp 1666464484
transform 1 0 9476 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_103
timestamp 1666464484
transform 1 0 10580 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_115
timestamp 1666464484
transform 1 0 11684 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_119
timestamp 1666464484
transform 1 0 12052 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_121
timestamp 1666464484
transform 1 0 12236 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_133
timestamp 1666464484
transform 1 0 13340 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_145
timestamp 1666464484
transform 1 0 14444 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_149
timestamp 1666464484
transform 1 0 14812 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_151
timestamp 1666464484
transform 1 0 14996 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_163
timestamp 1666464484
transform 1 0 16100 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_175
timestamp 1666464484
transform 1 0 17204 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_179
timestamp 1666464484
transform 1 0 17572 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1666464484
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1666464484
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_205
timestamp 1666464484
transform 1 0 19964 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_209
timestamp 1666464484
transform 1 0 20332 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_211
timestamp 1666464484
transform 1 0 20516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_223
timestamp 1666464484
transform 1 0 21620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_235
timestamp 1666464484
transform 1 0 22724 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_239
timestamp 1666464484
transform 1 0 23092 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_241
timestamp 1666464484
transform 1 0 23276 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_253
timestamp 1666464484
transform 1 0 24380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_265
timestamp 1666464484
transform 1 0 25484 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_269
timestamp 1666464484
transform 1 0 25852 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_271
timestamp 1666464484
transform 1 0 26036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_283
timestamp 1666464484
transform 1 0 27140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_295
timestamp 1666464484
transform 1 0 28244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_299
timestamp 1666464484
transform 1 0 28612 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_301
timestamp 1666464484
transform 1 0 28796 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_313
timestamp 1666464484
transform 1 0 29900 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_325
timestamp 1666464484
transform 1 0 31004 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_329
timestamp 1666464484
transform 1 0 31372 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_331
timestamp 1666464484
transform 1 0 31556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_343
timestamp 1666464484
transform 1 0 32660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_355
timestamp 1666464484
transform 1 0 33764 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_359
timestamp 1666464484
transform 1 0 34132 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1666464484
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1666464484
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_385
timestamp 1666464484
transform 1 0 36524 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_389
timestamp 1666464484
transform 1 0 36892 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_391
timestamp 1666464484
transform 1 0 37076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_403
timestamp 1666464484
transform 1 0 38180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_415
timestamp 1666464484
transform 1 0 39284 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_419
timestamp 1666464484
transform 1 0 39652 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_421
timestamp 1666464484
transform 1 0 39836 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_433
timestamp 1666464484
transform 1 0 40940 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_445
timestamp 1666464484
transform 1 0 42044 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_449
timestamp 1666464484
transform 1 0 42412 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_451
timestamp 1666464484
transform 1 0 42596 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_463
timestamp 1666464484
transform 1 0 43700 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_475
timestamp 1666464484
transform 1 0 44804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_479
timestamp 1666464484
transform 1 0 45172 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_481
timestamp 1666464484
transform 1 0 45356 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_493
timestamp 1666464484
transform 1 0 46460 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_505
timestamp 1666464484
transform 1 0 47564 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_509
timestamp 1666464484
transform 1 0 47932 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_511
timestamp 1666464484
transform 1 0 48116 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_523
timestamp 1666464484
transform 1 0 49220 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_535
timestamp 1666464484
transform 1 0 50324 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_539
timestamp 1666464484
transform 1 0 50692 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1666464484
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_553
timestamp 1666464484
transform 1 0 51980 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_565
timestamp 1666464484
transform 1 0 53084 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_569
timestamp 1666464484
transform 1 0 53452 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_571
timestamp 1666464484
transform 1 0 53636 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_583
timestamp 1666464484
transform 1 0 54740 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_595
timestamp 1666464484
transform 1 0 55844 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_599
timestamp 1666464484
transform 1 0 56212 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_601
timestamp 1666464484
transform 1 0 56396 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_613
timestamp 1666464484
transform 1 0 57500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_16
timestamp 1666464484
transform 1 0 2576 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_28
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_40
timestamp 1666464484
transform 1 0 4784 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_44
timestamp 1666464484
transform 1 0 5152 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_46
timestamp 1666464484
transform 1 0 5336 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_58
timestamp 1666464484
transform 1 0 6440 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_70
timestamp 1666464484
transform 1 0 7544 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_74
timestamp 1666464484
transform 1 0 7912 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_76
timestamp 1666464484
transform 1 0 8096 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_88
timestamp 1666464484
transform 1 0 9200 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_100
timestamp 1666464484
transform 1 0 10304 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_104
timestamp 1666464484
transform 1 0 10672 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_106
timestamp 1666464484
transform 1 0 10856 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_118
timestamp 1666464484
transform 1 0 11960 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_130
timestamp 1666464484
transform 1 0 13064 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_134
timestamp 1666464484
transform 1 0 13432 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_136
timestamp 1666464484
transform 1 0 13616 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_148
timestamp 1666464484
transform 1 0 14720 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_160
timestamp 1666464484
transform 1 0 15824 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_164
timestamp 1666464484
transform 1 0 16192 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_166
timestamp 1666464484
transform 1 0 16376 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_178
timestamp 1666464484
transform 1 0 17480 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_190
timestamp 1666464484
transform 1 0 18584 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_194
timestamp 1666464484
transform 1 0 18952 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_196
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_208
timestamp 1666464484
transform 1 0 20240 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_220
timestamp 1666464484
transform 1 0 21344 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_224
timestamp 1666464484
transform 1 0 21712 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_226
timestamp 1666464484
transform 1 0 21896 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_238
timestamp 1666464484
transform 1 0 23000 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_250
timestamp 1666464484
transform 1 0 24104 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_254
timestamp 1666464484
transform 1 0 24472 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_256
timestamp 1666464484
transform 1 0 24656 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_268
timestamp 1666464484
transform 1 0 25760 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_280
timestamp 1666464484
transform 1 0 26864 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_284
timestamp 1666464484
transform 1 0 27232 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_286
timestamp 1666464484
transform 1 0 27416 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_298
timestamp 1666464484
transform 1 0 28520 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_310
timestamp 1666464484
transform 1 0 29624 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_314
timestamp 1666464484
transform 1 0 29992 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_316
timestamp 1666464484
transform 1 0 30176 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_328
timestamp 1666464484
transform 1 0 31280 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_340
timestamp 1666464484
transform 1 0 32384 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_344
timestamp 1666464484
transform 1 0 32752 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_346
timestamp 1666464484
transform 1 0 32936 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_358
timestamp 1666464484
transform 1 0 34040 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_370
timestamp 1666464484
transform 1 0 35144 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_374
timestamp 1666464484
transform 1 0 35512 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_376
timestamp 1666464484
transform 1 0 35696 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_388
timestamp 1666464484
transform 1 0 36800 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_400
timestamp 1666464484
transform 1 0 37904 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_404
timestamp 1666464484
transform 1 0 38272 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_406
timestamp 1666464484
transform 1 0 38456 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_418
timestamp 1666464484
transform 1 0 39560 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_430
timestamp 1666464484
transform 1 0 40664 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_434
timestamp 1666464484
transform 1 0 41032 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_436
timestamp 1666464484
transform 1 0 41216 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_448
timestamp 1666464484
transform 1 0 42320 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_460
timestamp 1666464484
transform 1 0 43424 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_464
timestamp 1666464484
transform 1 0 43792 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_466
timestamp 1666464484
transform 1 0 43976 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_478
timestamp 1666464484
transform 1 0 45080 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_490
timestamp 1666464484
transform 1 0 46184 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_494
timestamp 1666464484
transform 1 0 46552 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_496
timestamp 1666464484
transform 1 0 46736 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_508
timestamp 1666464484
transform 1 0 47840 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_520
timestamp 1666464484
transform 1 0 48944 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_524
timestamp 1666464484
transform 1 0 49312 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_526
timestamp 1666464484
transform 1 0 49496 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_538
timestamp 1666464484
transform 1 0 50600 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_550
timestamp 1666464484
transform 1 0 51704 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_554
timestamp 1666464484
transform 1 0 52072 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_556
timestamp 1666464484
transform 1 0 52256 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_568
timestamp 1666464484
transform 1 0 53360 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_580
timestamp 1666464484
transform 1 0 54464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_584
timestamp 1666464484
transform 1 0 54832 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_586
timestamp 1666464484
transform 1 0 55016 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_598
timestamp 1666464484
transform 1 0 56120 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_610
timestamp 1666464484
transform 1 0 57224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_614
timestamp 1666464484
transform 1 0 57592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_616
timestamp 1666464484
transform 1 0 57776 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_624
timestamp 1666464484
transform 1 0 58512 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_31
timestamp 1666464484
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_43
timestamp 1666464484
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_55
timestamp 1666464484
transform 1 0 6164 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_59
timestamp 1666464484
transform 1 0 6532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_61
timestamp 1666464484
transform 1 0 6716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_73
timestamp 1666464484
transform 1 0 7820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_85
timestamp 1666464484
transform 1 0 8924 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_89
timestamp 1666464484
transform 1 0 9292 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_91
timestamp 1666464484
transform 1 0 9476 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_103
timestamp 1666464484
transform 1 0 10580 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_115
timestamp 1666464484
transform 1 0 11684 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_119
timestamp 1666464484
transform 1 0 12052 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_121
timestamp 1666464484
transform 1 0 12236 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_133
timestamp 1666464484
transform 1 0 13340 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_145
timestamp 1666464484
transform 1 0 14444 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_149
timestamp 1666464484
transform 1 0 14812 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_151
timestamp 1666464484
transform 1 0 14996 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_163
timestamp 1666464484
transform 1 0 16100 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_175
timestamp 1666464484
transform 1 0 17204 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_179
timestamp 1666464484
transform 1 0 17572 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1666464484
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1666464484
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_205
timestamp 1666464484
transform 1 0 19964 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_209
timestamp 1666464484
transform 1 0 20332 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_211
timestamp 1666464484
transform 1 0 20516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_223
timestamp 1666464484
transform 1 0 21620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_235
timestamp 1666464484
transform 1 0 22724 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_239
timestamp 1666464484
transform 1 0 23092 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_241
timestamp 1666464484
transform 1 0 23276 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_253
timestamp 1666464484
transform 1 0 24380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_265
timestamp 1666464484
transform 1 0 25484 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_269
timestamp 1666464484
transform 1 0 25852 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_271
timestamp 1666464484
transform 1 0 26036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_283
timestamp 1666464484
transform 1 0 27140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_295
timestamp 1666464484
transform 1 0 28244 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_299
timestamp 1666464484
transform 1 0 28612 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_301
timestamp 1666464484
transform 1 0 28796 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_313
timestamp 1666464484
transform 1 0 29900 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_325
timestamp 1666464484
transform 1 0 31004 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_329
timestamp 1666464484
transform 1 0 31372 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_331
timestamp 1666464484
transform 1 0 31556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_343
timestamp 1666464484
transform 1 0 32660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_355
timestamp 1666464484
transform 1 0 33764 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_359
timestamp 1666464484
transform 1 0 34132 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1666464484
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1666464484
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_385
timestamp 1666464484
transform 1 0 36524 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_389
timestamp 1666464484
transform 1 0 36892 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_391
timestamp 1666464484
transform 1 0 37076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_403
timestamp 1666464484
transform 1 0 38180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_415
timestamp 1666464484
transform 1 0 39284 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_419
timestamp 1666464484
transform 1 0 39652 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_421
timestamp 1666464484
transform 1 0 39836 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_433
timestamp 1666464484
transform 1 0 40940 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_445
timestamp 1666464484
transform 1 0 42044 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_449
timestamp 1666464484
transform 1 0 42412 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_451
timestamp 1666464484
transform 1 0 42596 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_463
timestamp 1666464484
transform 1 0 43700 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_475
timestamp 1666464484
transform 1 0 44804 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_479
timestamp 1666464484
transform 1 0 45172 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_481
timestamp 1666464484
transform 1 0 45356 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_493
timestamp 1666464484
transform 1 0 46460 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_505
timestamp 1666464484
transform 1 0 47564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_509
timestamp 1666464484
transform 1 0 47932 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_511
timestamp 1666464484
transform 1 0 48116 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_523
timestamp 1666464484
transform 1 0 49220 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_535
timestamp 1666464484
transform 1 0 50324 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_539
timestamp 1666464484
transform 1 0 50692 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1666464484
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_553
timestamp 1666464484
transform 1 0 51980 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_565
timestamp 1666464484
transform 1 0 53084 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_569
timestamp 1666464484
transform 1 0 53452 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_571
timestamp 1666464484
transform 1 0 53636 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_583
timestamp 1666464484
transform 1 0 54740 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_595
timestamp 1666464484
transform 1 0 55844 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_599
timestamp 1666464484
transform 1 0 56212 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_601
timestamp 1666464484
transform 1 0 56396 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_613
timestamp 1666464484
transform 1 0 57500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_16
timestamp 1666464484
transform 1 0 2576 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_28
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_40
timestamp 1666464484
transform 1 0 4784 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_44
timestamp 1666464484
transform 1 0 5152 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_46
timestamp 1666464484
transform 1 0 5336 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_58
timestamp 1666464484
transform 1 0 6440 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_70
timestamp 1666464484
transform 1 0 7544 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_74
timestamp 1666464484
transform 1 0 7912 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_76
timestamp 1666464484
transform 1 0 8096 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_88
timestamp 1666464484
transform 1 0 9200 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_100
timestamp 1666464484
transform 1 0 10304 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_104
timestamp 1666464484
transform 1 0 10672 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_106
timestamp 1666464484
transform 1 0 10856 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_118
timestamp 1666464484
transform 1 0 11960 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_130
timestamp 1666464484
transform 1 0 13064 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_134
timestamp 1666464484
transform 1 0 13432 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_136
timestamp 1666464484
transform 1 0 13616 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_148
timestamp 1666464484
transform 1 0 14720 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_160
timestamp 1666464484
transform 1 0 15824 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_164
timestamp 1666464484
transform 1 0 16192 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_166
timestamp 1666464484
transform 1 0 16376 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_178
timestamp 1666464484
transform 1 0 17480 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_190
timestamp 1666464484
transform 1 0 18584 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_194
timestamp 1666464484
transform 1 0 18952 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_196
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_208
timestamp 1666464484
transform 1 0 20240 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_220
timestamp 1666464484
transform 1 0 21344 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_224
timestamp 1666464484
transform 1 0 21712 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_226
timestamp 1666464484
transform 1 0 21896 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_238
timestamp 1666464484
transform 1 0 23000 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_250
timestamp 1666464484
transform 1 0 24104 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_254
timestamp 1666464484
transform 1 0 24472 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_256
timestamp 1666464484
transform 1 0 24656 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_268
timestamp 1666464484
transform 1 0 25760 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_280
timestamp 1666464484
transform 1 0 26864 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_284
timestamp 1666464484
transform 1 0 27232 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_286
timestamp 1666464484
transform 1 0 27416 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_298
timestamp 1666464484
transform 1 0 28520 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_310
timestamp 1666464484
transform 1 0 29624 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_314
timestamp 1666464484
transform 1 0 29992 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_316
timestamp 1666464484
transform 1 0 30176 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_328
timestamp 1666464484
transform 1 0 31280 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_340
timestamp 1666464484
transform 1 0 32384 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_344
timestamp 1666464484
transform 1 0 32752 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_346
timestamp 1666464484
transform 1 0 32936 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_358
timestamp 1666464484
transform 1 0 34040 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_370
timestamp 1666464484
transform 1 0 35144 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_374
timestamp 1666464484
transform 1 0 35512 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_376
timestamp 1666464484
transform 1 0 35696 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_388
timestamp 1666464484
transform 1 0 36800 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_400
timestamp 1666464484
transform 1 0 37904 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_404
timestamp 1666464484
transform 1 0 38272 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_406
timestamp 1666464484
transform 1 0 38456 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_418
timestamp 1666464484
transform 1 0 39560 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_430
timestamp 1666464484
transform 1 0 40664 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_434
timestamp 1666464484
transform 1 0 41032 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_436
timestamp 1666464484
transform 1 0 41216 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_448
timestamp 1666464484
transform 1 0 42320 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_460
timestamp 1666464484
transform 1 0 43424 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_464
timestamp 1666464484
transform 1 0 43792 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_466
timestamp 1666464484
transform 1 0 43976 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_478
timestamp 1666464484
transform 1 0 45080 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_490
timestamp 1666464484
transform 1 0 46184 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_494
timestamp 1666464484
transform 1 0 46552 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_496
timestamp 1666464484
transform 1 0 46736 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_508
timestamp 1666464484
transform 1 0 47840 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_520
timestamp 1666464484
transform 1 0 48944 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_524
timestamp 1666464484
transform 1 0 49312 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_526
timestamp 1666464484
transform 1 0 49496 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_538
timestamp 1666464484
transform 1 0 50600 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_550
timestamp 1666464484
transform 1 0 51704 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_554
timestamp 1666464484
transform 1 0 52072 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_556
timestamp 1666464484
transform 1 0 52256 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_568
timestamp 1666464484
transform 1 0 53360 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_580
timestamp 1666464484
transform 1 0 54464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_584
timestamp 1666464484
transform 1 0 54832 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_586
timestamp 1666464484
transform 1 0 55016 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_598
timestamp 1666464484
transform 1 0 56120 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_610
timestamp 1666464484
transform 1 0 57224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_614
timestamp 1666464484
transform 1 0 57592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_616
timestamp 1666464484
transform 1 0 57776 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_624
timestamp 1666464484
transform 1 0 58512 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666464484
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_27
timestamp 1666464484
transform 1 0 3588 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_31
timestamp 1666464484
transform 1 0 3956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_43
timestamp 1666464484
transform 1 0 5060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_55
timestamp 1666464484
transform 1 0 6164 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_59
timestamp 1666464484
transform 1 0 6532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_61
timestamp 1666464484
transform 1 0 6716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_73
timestamp 1666464484
transform 1 0 7820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_85
timestamp 1666464484
transform 1 0 8924 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_89
timestamp 1666464484
transform 1 0 9292 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_91
timestamp 1666464484
transform 1 0 9476 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_103
timestamp 1666464484
transform 1 0 10580 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_115
timestamp 1666464484
transform 1 0 11684 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_119
timestamp 1666464484
transform 1 0 12052 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_121
timestamp 1666464484
transform 1 0 12236 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_133
timestamp 1666464484
transform 1 0 13340 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_145
timestamp 1666464484
transform 1 0 14444 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_149
timestamp 1666464484
transform 1 0 14812 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_151
timestamp 1666464484
transform 1 0 14996 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_163
timestamp 1666464484
transform 1 0 16100 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_175
timestamp 1666464484
transform 1 0 17204 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_179
timestamp 1666464484
transform 1 0 17572 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1666464484
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1666464484
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_205
timestamp 1666464484
transform 1 0 19964 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_209
timestamp 1666464484
transform 1 0 20332 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_211
timestamp 1666464484
transform 1 0 20516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_223
timestamp 1666464484
transform 1 0 21620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_235
timestamp 1666464484
transform 1 0 22724 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_239
timestamp 1666464484
transform 1 0 23092 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_241
timestamp 1666464484
transform 1 0 23276 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_253
timestamp 1666464484
transform 1 0 24380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_265
timestamp 1666464484
transform 1 0 25484 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_269
timestamp 1666464484
transform 1 0 25852 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_271
timestamp 1666464484
transform 1 0 26036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_283
timestamp 1666464484
transform 1 0 27140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_295
timestamp 1666464484
transform 1 0 28244 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_299
timestamp 1666464484
transform 1 0 28612 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_301
timestamp 1666464484
transform 1 0 28796 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_313
timestamp 1666464484
transform 1 0 29900 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_325
timestamp 1666464484
transform 1 0 31004 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_329
timestamp 1666464484
transform 1 0 31372 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_331
timestamp 1666464484
transform 1 0 31556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_343
timestamp 1666464484
transform 1 0 32660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_355
timestamp 1666464484
transform 1 0 33764 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_359
timestamp 1666464484
transform 1 0 34132 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1666464484
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1666464484
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_385
timestamp 1666464484
transform 1 0 36524 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_389
timestamp 1666464484
transform 1 0 36892 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_391
timestamp 1666464484
transform 1 0 37076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_403
timestamp 1666464484
transform 1 0 38180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_415
timestamp 1666464484
transform 1 0 39284 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_419
timestamp 1666464484
transform 1 0 39652 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_421
timestamp 1666464484
transform 1 0 39836 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_433
timestamp 1666464484
transform 1 0 40940 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_445
timestamp 1666464484
transform 1 0 42044 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_449
timestamp 1666464484
transform 1 0 42412 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_451
timestamp 1666464484
transform 1 0 42596 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_463
timestamp 1666464484
transform 1 0 43700 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_475
timestamp 1666464484
transform 1 0 44804 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_479
timestamp 1666464484
transform 1 0 45172 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_481
timestamp 1666464484
transform 1 0 45356 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_493
timestamp 1666464484
transform 1 0 46460 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_505
timestamp 1666464484
transform 1 0 47564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_509
timestamp 1666464484
transform 1 0 47932 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_511
timestamp 1666464484
transform 1 0 48116 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_523
timestamp 1666464484
transform 1 0 49220 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_535
timestamp 1666464484
transform 1 0 50324 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_539
timestamp 1666464484
transform 1 0 50692 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1666464484
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_553
timestamp 1666464484
transform 1 0 51980 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_565
timestamp 1666464484
transform 1 0 53084 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_569
timestamp 1666464484
transform 1 0 53452 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_571
timestamp 1666464484
transform 1 0 53636 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_583
timestamp 1666464484
transform 1 0 54740 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_595
timestamp 1666464484
transform 1 0 55844 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_599
timestamp 1666464484
transform 1 0 56212 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_601
timestamp 1666464484
transform 1 0 56396 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_613
timestamp 1666464484
transform 1 0 57500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_16
timestamp 1666464484
transform 1 0 2576 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_28
timestamp 1666464484
transform 1 0 3680 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_40
timestamp 1666464484
transform 1 0 4784 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_44
timestamp 1666464484
transform 1 0 5152 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_46
timestamp 1666464484
transform 1 0 5336 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_58
timestamp 1666464484
transform 1 0 6440 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_70
timestamp 1666464484
transform 1 0 7544 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_74
timestamp 1666464484
transform 1 0 7912 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_76
timestamp 1666464484
transform 1 0 8096 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_88
timestamp 1666464484
transform 1 0 9200 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_100
timestamp 1666464484
transform 1 0 10304 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_104
timestamp 1666464484
transform 1 0 10672 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_106
timestamp 1666464484
transform 1 0 10856 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_118
timestamp 1666464484
transform 1 0 11960 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_130
timestamp 1666464484
transform 1 0 13064 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_134
timestamp 1666464484
transform 1 0 13432 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_136
timestamp 1666464484
transform 1 0 13616 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_148
timestamp 1666464484
transform 1 0 14720 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_160
timestamp 1666464484
transform 1 0 15824 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_164
timestamp 1666464484
transform 1 0 16192 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_166
timestamp 1666464484
transform 1 0 16376 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_178
timestamp 1666464484
transform 1 0 17480 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_190
timestamp 1666464484
transform 1 0 18584 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_194
timestamp 1666464484
transform 1 0 18952 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_196
timestamp 1666464484
transform 1 0 19136 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_208
timestamp 1666464484
transform 1 0 20240 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_220
timestamp 1666464484
transform 1 0 21344 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_224
timestamp 1666464484
transform 1 0 21712 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_226
timestamp 1666464484
transform 1 0 21896 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_238
timestamp 1666464484
transform 1 0 23000 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_250
timestamp 1666464484
transform 1 0 24104 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_254
timestamp 1666464484
transform 1 0 24472 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_256
timestamp 1666464484
transform 1 0 24656 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_268
timestamp 1666464484
transform 1 0 25760 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_280
timestamp 1666464484
transform 1 0 26864 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_284
timestamp 1666464484
transform 1 0 27232 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_286
timestamp 1666464484
transform 1 0 27416 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_298
timestamp 1666464484
transform 1 0 28520 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_310
timestamp 1666464484
transform 1 0 29624 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_314
timestamp 1666464484
transform 1 0 29992 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_316
timestamp 1666464484
transform 1 0 30176 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_328
timestamp 1666464484
transform 1 0 31280 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_340
timestamp 1666464484
transform 1 0 32384 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_344
timestamp 1666464484
transform 1 0 32752 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_346
timestamp 1666464484
transform 1 0 32936 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_358
timestamp 1666464484
transform 1 0 34040 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_370
timestamp 1666464484
transform 1 0 35144 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_374
timestamp 1666464484
transform 1 0 35512 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_376
timestamp 1666464484
transform 1 0 35696 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_388
timestamp 1666464484
transform 1 0 36800 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_400
timestamp 1666464484
transform 1 0 37904 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_404
timestamp 1666464484
transform 1 0 38272 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_406
timestamp 1666464484
transform 1 0 38456 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_418
timestamp 1666464484
transform 1 0 39560 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_430
timestamp 1666464484
transform 1 0 40664 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_434
timestamp 1666464484
transform 1 0 41032 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_436
timestamp 1666464484
transform 1 0 41216 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_448
timestamp 1666464484
transform 1 0 42320 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_460
timestamp 1666464484
transform 1 0 43424 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_464
timestamp 1666464484
transform 1 0 43792 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_466
timestamp 1666464484
transform 1 0 43976 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_478
timestamp 1666464484
transform 1 0 45080 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_490
timestamp 1666464484
transform 1 0 46184 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_494
timestamp 1666464484
transform 1 0 46552 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_496
timestamp 1666464484
transform 1 0 46736 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_508
timestamp 1666464484
transform 1 0 47840 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_520
timestamp 1666464484
transform 1 0 48944 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_524
timestamp 1666464484
transform 1 0 49312 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_526
timestamp 1666464484
transform 1 0 49496 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_538
timestamp 1666464484
transform 1 0 50600 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_550
timestamp 1666464484
transform 1 0 51704 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_554
timestamp 1666464484
transform 1 0 52072 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_556
timestamp 1666464484
transform 1 0 52256 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_568
timestamp 1666464484
transform 1 0 53360 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_580
timestamp 1666464484
transform 1 0 54464 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_584
timestamp 1666464484
transform 1 0 54832 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_586
timestamp 1666464484
transform 1 0 55016 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_598
timestamp 1666464484
transform 1 0 56120 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_610
timestamp 1666464484
transform 1 0 57224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_614
timestamp 1666464484
transform 1 0 57592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_616
timestamp 1666464484
transform 1 0 57776 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_624
timestamp 1666464484
transform 1 0 58512 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666464484
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_27
timestamp 1666464484
transform 1 0 3588 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_31
timestamp 1666464484
transform 1 0 3956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_43
timestamp 1666464484
transform 1 0 5060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_55
timestamp 1666464484
transform 1 0 6164 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_59
timestamp 1666464484
transform 1 0 6532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_61
timestamp 1666464484
transform 1 0 6716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_73
timestamp 1666464484
transform 1 0 7820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_85
timestamp 1666464484
transform 1 0 8924 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_89
timestamp 1666464484
transform 1 0 9292 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_91
timestamp 1666464484
transform 1 0 9476 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_103
timestamp 1666464484
transform 1 0 10580 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_115
timestamp 1666464484
transform 1 0 11684 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_119
timestamp 1666464484
transform 1 0 12052 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_121
timestamp 1666464484
transform 1 0 12236 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_133
timestamp 1666464484
transform 1 0 13340 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_145
timestamp 1666464484
transform 1 0 14444 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_149
timestamp 1666464484
transform 1 0 14812 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_151
timestamp 1666464484
transform 1 0 14996 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_163
timestamp 1666464484
transform 1 0 16100 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_175
timestamp 1666464484
transform 1 0 17204 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_179
timestamp 1666464484
transform 1 0 17572 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1666464484
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1666464484
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_205
timestamp 1666464484
transform 1 0 19964 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_209
timestamp 1666464484
transform 1 0 20332 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_211
timestamp 1666464484
transform 1 0 20516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_223
timestamp 1666464484
transform 1 0 21620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_235
timestamp 1666464484
transform 1 0 22724 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_239
timestamp 1666464484
transform 1 0 23092 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_241
timestamp 1666464484
transform 1 0 23276 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_253
timestamp 1666464484
transform 1 0 24380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_265
timestamp 1666464484
transform 1 0 25484 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_269
timestamp 1666464484
transform 1 0 25852 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_271
timestamp 1666464484
transform 1 0 26036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_283
timestamp 1666464484
transform 1 0 27140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_295
timestamp 1666464484
transform 1 0 28244 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_299
timestamp 1666464484
transform 1 0 28612 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_301
timestamp 1666464484
transform 1 0 28796 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_313
timestamp 1666464484
transform 1 0 29900 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_325
timestamp 1666464484
transform 1 0 31004 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_329
timestamp 1666464484
transform 1 0 31372 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_331
timestamp 1666464484
transform 1 0 31556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_343
timestamp 1666464484
transform 1 0 32660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_355
timestamp 1666464484
transform 1 0 33764 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_359
timestamp 1666464484
transform 1 0 34132 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1666464484
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1666464484
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_385
timestamp 1666464484
transform 1 0 36524 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_389
timestamp 1666464484
transform 1 0 36892 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_391
timestamp 1666464484
transform 1 0 37076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_403
timestamp 1666464484
transform 1 0 38180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_415
timestamp 1666464484
transform 1 0 39284 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_419
timestamp 1666464484
transform 1 0 39652 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_421
timestamp 1666464484
transform 1 0 39836 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_433
timestamp 1666464484
transform 1 0 40940 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_445
timestamp 1666464484
transform 1 0 42044 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_449
timestamp 1666464484
transform 1 0 42412 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_451
timestamp 1666464484
transform 1 0 42596 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_463
timestamp 1666464484
transform 1 0 43700 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_475
timestamp 1666464484
transform 1 0 44804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_479
timestamp 1666464484
transform 1 0 45172 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_481
timestamp 1666464484
transform 1 0 45356 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_493
timestamp 1666464484
transform 1 0 46460 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_505
timestamp 1666464484
transform 1 0 47564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_509
timestamp 1666464484
transform 1 0 47932 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_511
timestamp 1666464484
transform 1 0 48116 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_523
timestamp 1666464484
transform 1 0 49220 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_535
timestamp 1666464484
transform 1 0 50324 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_539
timestamp 1666464484
transform 1 0 50692 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1666464484
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_553
timestamp 1666464484
transform 1 0 51980 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_565
timestamp 1666464484
transform 1 0 53084 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_569
timestamp 1666464484
transform 1 0 53452 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_571
timestamp 1666464484
transform 1 0 53636 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_583
timestamp 1666464484
transform 1 0 54740 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_595
timestamp 1666464484
transform 1 0 55844 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_599
timestamp 1666464484
transform 1 0 56212 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_601
timestamp 1666464484
transform 1 0 56396 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_613
timestamp 1666464484
transform 1 0 57500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_16
timestamp 1666464484
transform 1 0 2576 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_28
timestamp 1666464484
transform 1 0 3680 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_40
timestamp 1666464484
transform 1 0 4784 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_44
timestamp 1666464484
transform 1 0 5152 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_46
timestamp 1666464484
transform 1 0 5336 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_58
timestamp 1666464484
transform 1 0 6440 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_70
timestamp 1666464484
transform 1 0 7544 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_74
timestamp 1666464484
transform 1 0 7912 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_76
timestamp 1666464484
transform 1 0 8096 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_88
timestamp 1666464484
transform 1 0 9200 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_100
timestamp 1666464484
transform 1 0 10304 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_104
timestamp 1666464484
transform 1 0 10672 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_106
timestamp 1666464484
transform 1 0 10856 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_118
timestamp 1666464484
transform 1 0 11960 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_130
timestamp 1666464484
transform 1 0 13064 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_134
timestamp 1666464484
transform 1 0 13432 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_136
timestamp 1666464484
transform 1 0 13616 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_148
timestamp 1666464484
transform 1 0 14720 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_160
timestamp 1666464484
transform 1 0 15824 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_164
timestamp 1666464484
transform 1 0 16192 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_166
timestamp 1666464484
transform 1 0 16376 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_178
timestamp 1666464484
transform 1 0 17480 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_190
timestamp 1666464484
transform 1 0 18584 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_194
timestamp 1666464484
transform 1 0 18952 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_196
timestamp 1666464484
transform 1 0 19136 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_208
timestamp 1666464484
transform 1 0 20240 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_220
timestamp 1666464484
transform 1 0 21344 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_224
timestamp 1666464484
transform 1 0 21712 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_226
timestamp 1666464484
transform 1 0 21896 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_238
timestamp 1666464484
transform 1 0 23000 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_250
timestamp 1666464484
transform 1 0 24104 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_254
timestamp 1666464484
transform 1 0 24472 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_256
timestamp 1666464484
transform 1 0 24656 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_268
timestamp 1666464484
transform 1 0 25760 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_280
timestamp 1666464484
transform 1 0 26864 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_284
timestamp 1666464484
transform 1 0 27232 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_286
timestamp 1666464484
transform 1 0 27416 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_298
timestamp 1666464484
transform 1 0 28520 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_310
timestamp 1666464484
transform 1 0 29624 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_314
timestamp 1666464484
transform 1 0 29992 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_316
timestamp 1666464484
transform 1 0 30176 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_328
timestamp 1666464484
transform 1 0 31280 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_340
timestamp 1666464484
transform 1 0 32384 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_344
timestamp 1666464484
transform 1 0 32752 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_346
timestamp 1666464484
transform 1 0 32936 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_358
timestamp 1666464484
transform 1 0 34040 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_370
timestamp 1666464484
transform 1 0 35144 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_374
timestamp 1666464484
transform 1 0 35512 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_376
timestamp 1666464484
transform 1 0 35696 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_388
timestamp 1666464484
transform 1 0 36800 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_400
timestamp 1666464484
transform 1 0 37904 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_404
timestamp 1666464484
transform 1 0 38272 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_406
timestamp 1666464484
transform 1 0 38456 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_418
timestamp 1666464484
transform 1 0 39560 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_430
timestamp 1666464484
transform 1 0 40664 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_434
timestamp 1666464484
transform 1 0 41032 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_436
timestamp 1666464484
transform 1 0 41216 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_448
timestamp 1666464484
transform 1 0 42320 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_460
timestamp 1666464484
transform 1 0 43424 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_464
timestamp 1666464484
transform 1 0 43792 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_466
timestamp 1666464484
transform 1 0 43976 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_478
timestamp 1666464484
transform 1 0 45080 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_490
timestamp 1666464484
transform 1 0 46184 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_494
timestamp 1666464484
transform 1 0 46552 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_496
timestamp 1666464484
transform 1 0 46736 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_508
timestamp 1666464484
transform 1 0 47840 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_520
timestamp 1666464484
transform 1 0 48944 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_524
timestamp 1666464484
transform 1 0 49312 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_526
timestamp 1666464484
transform 1 0 49496 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_538
timestamp 1666464484
transform 1 0 50600 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_550
timestamp 1666464484
transform 1 0 51704 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_554
timestamp 1666464484
transform 1 0 52072 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_556
timestamp 1666464484
transform 1 0 52256 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_568
timestamp 1666464484
transform 1 0 53360 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_580
timestamp 1666464484
transform 1 0 54464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_584
timestamp 1666464484
transform 1 0 54832 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_586
timestamp 1666464484
transform 1 0 55016 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_598
timestamp 1666464484
transform 1 0 56120 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_610
timestamp 1666464484
transform 1 0 57224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_614
timestamp 1666464484
transform 1 0 57592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_616
timestamp 1666464484
transform 1 0 57776 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_624
timestamp 1666464484
transform 1 0 58512 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666464484
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_27
timestamp 1666464484
transform 1 0 3588 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_31
timestamp 1666464484
transform 1 0 3956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_43
timestamp 1666464484
transform 1 0 5060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_55
timestamp 1666464484
transform 1 0 6164 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_59
timestamp 1666464484
transform 1 0 6532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_61
timestamp 1666464484
transform 1 0 6716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_73
timestamp 1666464484
transform 1 0 7820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_85
timestamp 1666464484
transform 1 0 8924 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_89
timestamp 1666464484
transform 1 0 9292 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_91
timestamp 1666464484
transform 1 0 9476 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_103
timestamp 1666464484
transform 1 0 10580 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_115
timestamp 1666464484
transform 1 0 11684 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_119
timestamp 1666464484
transform 1 0 12052 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_121
timestamp 1666464484
transform 1 0 12236 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_133
timestamp 1666464484
transform 1 0 13340 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_145
timestamp 1666464484
transform 1 0 14444 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_149
timestamp 1666464484
transform 1 0 14812 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_151
timestamp 1666464484
transform 1 0 14996 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_163
timestamp 1666464484
transform 1 0 16100 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_175
timestamp 1666464484
transform 1 0 17204 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_179
timestamp 1666464484
transform 1 0 17572 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1666464484
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1666464484
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_205
timestamp 1666464484
transform 1 0 19964 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_209
timestamp 1666464484
transform 1 0 20332 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_211
timestamp 1666464484
transform 1 0 20516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_223
timestamp 1666464484
transform 1 0 21620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_235
timestamp 1666464484
transform 1 0 22724 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_239
timestamp 1666464484
transform 1 0 23092 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_241
timestamp 1666464484
transform 1 0 23276 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_253
timestamp 1666464484
transform 1 0 24380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_265
timestamp 1666464484
transform 1 0 25484 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_269
timestamp 1666464484
transform 1 0 25852 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_271
timestamp 1666464484
transform 1 0 26036 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_283
timestamp 1666464484
transform 1 0 27140 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_295
timestamp 1666464484
transform 1 0 28244 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_299
timestamp 1666464484
transform 1 0 28612 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_301
timestamp 1666464484
transform 1 0 28796 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_313
timestamp 1666464484
transform 1 0 29900 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_325
timestamp 1666464484
transform 1 0 31004 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_329
timestamp 1666464484
transform 1 0 31372 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_331
timestamp 1666464484
transform 1 0 31556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_343
timestamp 1666464484
transform 1 0 32660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_355
timestamp 1666464484
transform 1 0 33764 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_359
timestamp 1666464484
transform 1 0 34132 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1666464484
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1666464484
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_385
timestamp 1666464484
transform 1 0 36524 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_389
timestamp 1666464484
transform 1 0 36892 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_391
timestamp 1666464484
transform 1 0 37076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_403
timestamp 1666464484
transform 1 0 38180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_415
timestamp 1666464484
transform 1 0 39284 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_419
timestamp 1666464484
transform 1 0 39652 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_421
timestamp 1666464484
transform 1 0 39836 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_433
timestamp 1666464484
transform 1 0 40940 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_445
timestamp 1666464484
transform 1 0 42044 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_449
timestamp 1666464484
transform 1 0 42412 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_451
timestamp 1666464484
transform 1 0 42596 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_463
timestamp 1666464484
transform 1 0 43700 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_475
timestamp 1666464484
transform 1 0 44804 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_479
timestamp 1666464484
transform 1 0 45172 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_481
timestamp 1666464484
transform 1 0 45356 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_493
timestamp 1666464484
transform 1 0 46460 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_505
timestamp 1666464484
transform 1 0 47564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_509
timestamp 1666464484
transform 1 0 47932 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_511
timestamp 1666464484
transform 1 0 48116 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_523
timestamp 1666464484
transform 1 0 49220 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_535
timestamp 1666464484
transform 1 0 50324 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_539
timestamp 1666464484
transform 1 0 50692 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1666464484
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_553
timestamp 1666464484
transform 1 0 51980 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_565
timestamp 1666464484
transform 1 0 53084 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_569
timestamp 1666464484
transform 1 0 53452 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_571
timestamp 1666464484
transform 1 0 53636 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_583
timestamp 1666464484
transform 1 0 54740 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_595
timestamp 1666464484
transform 1 0 55844 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_599
timestamp 1666464484
transform 1 0 56212 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_601
timestamp 1666464484
transform 1 0 56396 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_613
timestamp 1666464484
transform 1 0 57500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_16
timestamp 1666464484
transform 1 0 2576 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_28
timestamp 1666464484
transform 1 0 3680 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_40
timestamp 1666464484
transform 1 0 4784 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_44
timestamp 1666464484
transform 1 0 5152 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_46
timestamp 1666464484
transform 1 0 5336 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_58
timestamp 1666464484
transform 1 0 6440 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_70
timestamp 1666464484
transform 1 0 7544 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_74
timestamp 1666464484
transform 1 0 7912 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_76
timestamp 1666464484
transform 1 0 8096 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_88
timestamp 1666464484
transform 1 0 9200 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_100
timestamp 1666464484
transform 1 0 10304 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_104
timestamp 1666464484
transform 1 0 10672 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_106
timestamp 1666464484
transform 1 0 10856 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_118
timestamp 1666464484
transform 1 0 11960 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_130
timestamp 1666464484
transform 1 0 13064 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_134
timestamp 1666464484
transform 1 0 13432 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_136
timestamp 1666464484
transform 1 0 13616 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_148
timestamp 1666464484
transform 1 0 14720 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_160
timestamp 1666464484
transform 1 0 15824 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_164
timestamp 1666464484
transform 1 0 16192 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_166
timestamp 1666464484
transform 1 0 16376 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_178
timestamp 1666464484
transform 1 0 17480 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_190
timestamp 1666464484
transform 1 0 18584 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_194
timestamp 1666464484
transform 1 0 18952 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_196
timestamp 1666464484
transform 1 0 19136 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_208
timestamp 1666464484
transform 1 0 20240 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_220
timestamp 1666464484
transform 1 0 21344 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_224
timestamp 1666464484
transform 1 0 21712 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_226
timestamp 1666464484
transform 1 0 21896 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_238
timestamp 1666464484
transform 1 0 23000 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_250
timestamp 1666464484
transform 1 0 24104 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_254
timestamp 1666464484
transform 1 0 24472 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_256
timestamp 1666464484
transform 1 0 24656 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_268
timestamp 1666464484
transform 1 0 25760 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_280
timestamp 1666464484
transform 1 0 26864 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_284
timestamp 1666464484
transform 1 0 27232 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_286
timestamp 1666464484
transform 1 0 27416 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_298
timestamp 1666464484
transform 1 0 28520 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_310
timestamp 1666464484
transform 1 0 29624 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_314
timestamp 1666464484
transform 1 0 29992 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_316
timestamp 1666464484
transform 1 0 30176 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_328
timestamp 1666464484
transform 1 0 31280 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_340
timestamp 1666464484
transform 1 0 32384 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_344
timestamp 1666464484
transform 1 0 32752 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_346
timestamp 1666464484
transform 1 0 32936 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_358
timestamp 1666464484
transform 1 0 34040 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_370
timestamp 1666464484
transform 1 0 35144 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_374
timestamp 1666464484
transform 1 0 35512 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_376
timestamp 1666464484
transform 1 0 35696 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_388
timestamp 1666464484
transform 1 0 36800 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_400
timestamp 1666464484
transform 1 0 37904 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_404
timestamp 1666464484
transform 1 0 38272 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_406
timestamp 1666464484
transform 1 0 38456 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_418
timestamp 1666464484
transform 1 0 39560 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_430
timestamp 1666464484
transform 1 0 40664 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_434
timestamp 1666464484
transform 1 0 41032 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_436
timestamp 1666464484
transform 1 0 41216 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_448
timestamp 1666464484
transform 1 0 42320 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_460
timestamp 1666464484
transform 1 0 43424 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_464
timestamp 1666464484
transform 1 0 43792 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_466
timestamp 1666464484
transform 1 0 43976 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_478
timestamp 1666464484
transform 1 0 45080 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_490
timestamp 1666464484
transform 1 0 46184 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_494
timestamp 1666464484
transform 1 0 46552 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_496
timestamp 1666464484
transform 1 0 46736 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_508
timestamp 1666464484
transform 1 0 47840 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_520
timestamp 1666464484
transform 1 0 48944 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_524
timestamp 1666464484
transform 1 0 49312 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_526
timestamp 1666464484
transform 1 0 49496 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_538
timestamp 1666464484
transform 1 0 50600 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_550
timestamp 1666464484
transform 1 0 51704 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_554
timestamp 1666464484
transform 1 0 52072 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_556
timestamp 1666464484
transform 1 0 52256 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_568
timestamp 1666464484
transform 1 0 53360 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_580
timestamp 1666464484
transform 1 0 54464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_584
timestamp 1666464484
transform 1 0 54832 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_586
timestamp 1666464484
transform 1 0 55016 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_598
timestamp 1666464484
transform 1 0 56120 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_610
timestamp 1666464484
transform 1 0 57224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_614
timestamp 1666464484
transform 1 0 57592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_616
timestamp 1666464484
transform 1 0 57776 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_624
timestamp 1666464484
transform 1 0 58512 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666464484
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_27
timestamp 1666464484
transform 1 0 3588 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_31
timestamp 1666464484
transform 1 0 3956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_43
timestamp 1666464484
transform 1 0 5060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_55
timestamp 1666464484
transform 1 0 6164 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_59
timestamp 1666464484
transform 1 0 6532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_61
timestamp 1666464484
transform 1 0 6716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_73
timestamp 1666464484
transform 1 0 7820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_85
timestamp 1666464484
transform 1 0 8924 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_89
timestamp 1666464484
transform 1 0 9292 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_91
timestamp 1666464484
transform 1 0 9476 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_103
timestamp 1666464484
transform 1 0 10580 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_115
timestamp 1666464484
transform 1 0 11684 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_119
timestamp 1666464484
transform 1 0 12052 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_121
timestamp 1666464484
transform 1 0 12236 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_133
timestamp 1666464484
transform 1 0 13340 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_145
timestamp 1666464484
transform 1 0 14444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_149
timestamp 1666464484
transform 1 0 14812 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_151
timestamp 1666464484
transform 1 0 14996 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_163
timestamp 1666464484
transform 1 0 16100 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_175
timestamp 1666464484
transform 1 0 17204 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_179
timestamp 1666464484
transform 1 0 17572 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1666464484
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1666464484
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_205
timestamp 1666464484
transform 1 0 19964 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_209
timestamp 1666464484
transform 1 0 20332 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_211
timestamp 1666464484
transform 1 0 20516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_223
timestamp 1666464484
transform 1 0 21620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_235
timestamp 1666464484
transform 1 0 22724 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_239
timestamp 1666464484
transform 1 0 23092 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_241
timestamp 1666464484
transform 1 0 23276 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_253
timestamp 1666464484
transform 1 0 24380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_265
timestamp 1666464484
transform 1 0 25484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_269
timestamp 1666464484
transform 1 0 25852 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_271
timestamp 1666464484
transform 1 0 26036 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_283
timestamp 1666464484
transform 1 0 27140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_295
timestamp 1666464484
transform 1 0 28244 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_299
timestamp 1666464484
transform 1 0 28612 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_301
timestamp 1666464484
transform 1 0 28796 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_313
timestamp 1666464484
transform 1 0 29900 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_325
timestamp 1666464484
transform 1 0 31004 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_329
timestamp 1666464484
transform 1 0 31372 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_331
timestamp 1666464484
transform 1 0 31556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_343
timestamp 1666464484
transform 1 0 32660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_355
timestamp 1666464484
transform 1 0 33764 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_359
timestamp 1666464484
transform 1 0 34132 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1666464484
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1666464484
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_385
timestamp 1666464484
transform 1 0 36524 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_389
timestamp 1666464484
transform 1 0 36892 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_391
timestamp 1666464484
transform 1 0 37076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_403
timestamp 1666464484
transform 1 0 38180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_415
timestamp 1666464484
transform 1 0 39284 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_419
timestamp 1666464484
transform 1 0 39652 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_421
timestamp 1666464484
transform 1 0 39836 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_433
timestamp 1666464484
transform 1 0 40940 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_445
timestamp 1666464484
transform 1 0 42044 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_449
timestamp 1666464484
transform 1 0 42412 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_451
timestamp 1666464484
transform 1 0 42596 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_463
timestamp 1666464484
transform 1 0 43700 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_475
timestamp 1666464484
transform 1 0 44804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_479
timestamp 1666464484
transform 1 0 45172 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_481
timestamp 1666464484
transform 1 0 45356 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_493
timestamp 1666464484
transform 1 0 46460 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_505
timestamp 1666464484
transform 1 0 47564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_509
timestamp 1666464484
transform 1 0 47932 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_511
timestamp 1666464484
transform 1 0 48116 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_523
timestamp 1666464484
transform 1 0 49220 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_535
timestamp 1666464484
transform 1 0 50324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_539
timestamp 1666464484
transform 1 0 50692 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1666464484
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_553
timestamp 1666464484
transform 1 0 51980 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_565
timestamp 1666464484
transform 1 0 53084 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_569
timestamp 1666464484
transform 1 0 53452 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_571
timestamp 1666464484
transform 1 0 53636 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_583
timestamp 1666464484
transform 1 0 54740 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_595
timestamp 1666464484
transform 1 0 55844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_599
timestamp 1666464484
transform 1 0 56212 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_601
timestamp 1666464484
transform 1 0 56396 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_613
timestamp 1666464484
transform 1 0 57500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_16
timestamp 1666464484
transform 1 0 2576 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_28
timestamp 1666464484
transform 1 0 3680 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_40
timestamp 1666464484
transform 1 0 4784 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_44
timestamp 1666464484
transform 1 0 5152 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_46
timestamp 1666464484
transform 1 0 5336 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_58
timestamp 1666464484
transform 1 0 6440 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_70
timestamp 1666464484
transform 1 0 7544 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_74
timestamp 1666464484
transform 1 0 7912 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_76
timestamp 1666464484
transform 1 0 8096 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_88
timestamp 1666464484
transform 1 0 9200 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_100
timestamp 1666464484
transform 1 0 10304 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_104
timestamp 1666464484
transform 1 0 10672 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_106
timestamp 1666464484
transform 1 0 10856 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_118
timestamp 1666464484
transform 1 0 11960 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_130
timestamp 1666464484
transform 1 0 13064 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_134
timestamp 1666464484
transform 1 0 13432 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_136
timestamp 1666464484
transform 1 0 13616 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_148
timestamp 1666464484
transform 1 0 14720 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_160
timestamp 1666464484
transform 1 0 15824 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_164
timestamp 1666464484
transform 1 0 16192 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_166
timestamp 1666464484
transform 1 0 16376 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_178
timestamp 1666464484
transform 1 0 17480 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_190
timestamp 1666464484
transform 1 0 18584 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_194
timestamp 1666464484
transform 1 0 18952 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_196
timestamp 1666464484
transform 1 0 19136 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_208
timestamp 1666464484
transform 1 0 20240 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_220
timestamp 1666464484
transform 1 0 21344 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_224
timestamp 1666464484
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_226
timestamp 1666464484
transform 1 0 21896 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_238
timestamp 1666464484
transform 1 0 23000 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_250
timestamp 1666464484
transform 1 0 24104 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_254
timestamp 1666464484
transform 1 0 24472 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_256
timestamp 1666464484
transform 1 0 24656 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_268
timestamp 1666464484
transform 1 0 25760 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_280
timestamp 1666464484
transform 1 0 26864 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_284
timestamp 1666464484
transform 1 0 27232 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_286
timestamp 1666464484
transform 1 0 27416 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_298
timestamp 1666464484
transform 1 0 28520 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_310
timestamp 1666464484
transform 1 0 29624 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_314
timestamp 1666464484
transform 1 0 29992 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_316
timestamp 1666464484
transform 1 0 30176 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_328
timestamp 1666464484
transform 1 0 31280 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_340
timestamp 1666464484
transform 1 0 32384 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_344
timestamp 1666464484
transform 1 0 32752 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_346
timestamp 1666464484
transform 1 0 32936 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_358
timestamp 1666464484
transform 1 0 34040 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_370
timestamp 1666464484
transform 1 0 35144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_374
timestamp 1666464484
transform 1 0 35512 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_376
timestamp 1666464484
transform 1 0 35696 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_388
timestamp 1666464484
transform 1 0 36800 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_400
timestamp 1666464484
transform 1 0 37904 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_404
timestamp 1666464484
transform 1 0 38272 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_406
timestamp 1666464484
transform 1 0 38456 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_418
timestamp 1666464484
transform 1 0 39560 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_430
timestamp 1666464484
transform 1 0 40664 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_434
timestamp 1666464484
transform 1 0 41032 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_436
timestamp 1666464484
transform 1 0 41216 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_448
timestamp 1666464484
transform 1 0 42320 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_460
timestamp 1666464484
transform 1 0 43424 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_464
timestamp 1666464484
transform 1 0 43792 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_466
timestamp 1666464484
transform 1 0 43976 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_478
timestamp 1666464484
transform 1 0 45080 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_490
timestamp 1666464484
transform 1 0 46184 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_494
timestamp 1666464484
transform 1 0 46552 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_496
timestamp 1666464484
transform 1 0 46736 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_508
timestamp 1666464484
transform 1 0 47840 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_520
timestamp 1666464484
transform 1 0 48944 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_524
timestamp 1666464484
transform 1 0 49312 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_526
timestamp 1666464484
transform 1 0 49496 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_538
timestamp 1666464484
transform 1 0 50600 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_550
timestamp 1666464484
transform 1 0 51704 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_554
timestamp 1666464484
transform 1 0 52072 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_556
timestamp 1666464484
transform 1 0 52256 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_568
timestamp 1666464484
transform 1 0 53360 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_580
timestamp 1666464484
transform 1 0 54464 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_584
timestamp 1666464484
transform 1 0 54832 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_586
timestamp 1666464484
transform 1 0 55016 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_598
timestamp 1666464484
transform 1 0 56120 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_610
timestamp 1666464484
transform 1 0 57224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_614
timestamp 1666464484
transform 1 0 57592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_616
timestamp 1666464484
transform 1 0 57776 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_624
timestamp 1666464484
transform 1 0 58512 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1666464484
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1666464484
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_27
timestamp 1666464484
transform 1 0 3588 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_31
timestamp 1666464484
transform 1 0 3956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_43
timestamp 1666464484
transform 1 0 5060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_55
timestamp 1666464484
transform 1 0 6164 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_59
timestamp 1666464484
transform 1 0 6532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_61
timestamp 1666464484
transform 1 0 6716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_73
timestamp 1666464484
transform 1 0 7820 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_85
timestamp 1666464484
transform 1 0 8924 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_89
timestamp 1666464484
transform 1 0 9292 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_91
timestamp 1666464484
transform 1 0 9476 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_103
timestamp 1666464484
transform 1 0 10580 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_115
timestamp 1666464484
transform 1 0 11684 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_119
timestamp 1666464484
transform 1 0 12052 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_121
timestamp 1666464484
transform 1 0 12236 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_133
timestamp 1666464484
transform 1 0 13340 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_145
timestamp 1666464484
transform 1 0 14444 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_149
timestamp 1666464484
transform 1 0 14812 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_151
timestamp 1666464484
transform 1 0 14996 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_163
timestamp 1666464484
transform 1 0 16100 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_175
timestamp 1666464484
transform 1 0 17204 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_179
timestamp 1666464484
transform 1 0 17572 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1666464484
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1666464484
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_205
timestamp 1666464484
transform 1 0 19964 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_209
timestamp 1666464484
transform 1 0 20332 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_211
timestamp 1666464484
transform 1 0 20516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_223
timestamp 1666464484
transform 1 0 21620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_235
timestamp 1666464484
transform 1 0 22724 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_239
timestamp 1666464484
transform 1 0 23092 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_241
timestamp 1666464484
transform 1 0 23276 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_253
timestamp 1666464484
transform 1 0 24380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_265
timestamp 1666464484
transform 1 0 25484 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_269
timestamp 1666464484
transform 1 0 25852 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_271
timestamp 1666464484
transform 1 0 26036 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_283
timestamp 1666464484
transform 1 0 27140 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_295
timestamp 1666464484
transform 1 0 28244 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_299
timestamp 1666464484
transform 1 0 28612 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_301
timestamp 1666464484
transform 1 0 28796 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_313
timestamp 1666464484
transform 1 0 29900 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_325
timestamp 1666464484
transform 1 0 31004 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_329
timestamp 1666464484
transform 1 0 31372 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_331
timestamp 1666464484
transform 1 0 31556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_343
timestamp 1666464484
transform 1 0 32660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_355
timestamp 1666464484
transform 1 0 33764 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_359
timestamp 1666464484
transform 1 0 34132 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1666464484
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1666464484
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_385
timestamp 1666464484
transform 1 0 36524 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_389
timestamp 1666464484
transform 1 0 36892 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_391
timestamp 1666464484
transform 1 0 37076 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_403
timestamp 1666464484
transform 1 0 38180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_415
timestamp 1666464484
transform 1 0 39284 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_419
timestamp 1666464484
transform 1 0 39652 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_421
timestamp 1666464484
transform 1 0 39836 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_433
timestamp 1666464484
transform 1 0 40940 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_445
timestamp 1666464484
transform 1 0 42044 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_449
timestamp 1666464484
transform 1 0 42412 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_451
timestamp 1666464484
transform 1 0 42596 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_463
timestamp 1666464484
transform 1 0 43700 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_475
timestamp 1666464484
transform 1 0 44804 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_479
timestamp 1666464484
transform 1 0 45172 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_481
timestamp 1666464484
transform 1 0 45356 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_493
timestamp 1666464484
transform 1 0 46460 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_505
timestamp 1666464484
transform 1 0 47564 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_509
timestamp 1666464484
transform 1 0 47932 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_511
timestamp 1666464484
transform 1 0 48116 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_523
timestamp 1666464484
transform 1 0 49220 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_535
timestamp 1666464484
transform 1 0 50324 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_539
timestamp 1666464484
transform 1 0 50692 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1666464484
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_553
timestamp 1666464484
transform 1 0 51980 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_565
timestamp 1666464484
transform 1 0 53084 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_569
timestamp 1666464484
transform 1 0 53452 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_571
timestamp 1666464484
transform 1 0 53636 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_583
timestamp 1666464484
transform 1 0 54740 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_595
timestamp 1666464484
transform 1 0 55844 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_599
timestamp 1666464484
transform 1 0 56212 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_601
timestamp 1666464484
transform 1 0 56396 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_613
timestamp 1666464484
transform 1 0 57500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1666464484
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_16
timestamp 1666464484
transform 1 0 2576 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_28
timestamp 1666464484
transform 1 0 3680 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_40
timestamp 1666464484
transform 1 0 4784 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_44
timestamp 1666464484
transform 1 0 5152 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_46
timestamp 1666464484
transform 1 0 5336 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_58
timestamp 1666464484
transform 1 0 6440 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_70
timestamp 1666464484
transform 1 0 7544 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_74
timestamp 1666464484
transform 1 0 7912 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_76
timestamp 1666464484
transform 1 0 8096 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_88
timestamp 1666464484
transform 1 0 9200 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_100
timestamp 1666464484
transform 1 0 10304 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_104
timestamp 1666464484
transform 1 0 10672 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_106
timestamp 1666464484
transform 1 0 10856 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_118
timestamp 1666464484
transform 1 0 11960 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_130
timestamp 1666464484
transform 1 0 13064 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_134
timestamp 1666464484
transform 1 0 13432 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_136
timestamp 1666464484
transform 1 0 13616 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_148
timestamp 1666464484
transform 1 0 14720 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_160
timestamp 1666464484
transform 1 0 15824 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_164
timestamp 1666464484
transform 1 0 16192 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_166
timestamp 1666464484
transform 1 0 16376 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_178
timestamp 1666464484
transform 1 0 17480 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_190
timestamp 1666464484
transform 1 0 18584 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_194
timestamp 1666464484
transform 1 0 18952 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_196
timestamp 1666464484
transform 1 0 19136 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_208
timestamp 1666464484
transform 1 0 20240 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_220
timestamp 1666464484
transform 1 0 21344 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_224
timestamp 1666464484
transform 1 0 21712 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_226
timestamp 1666464484
transform 1 0 21896 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_238
timestamp 1666464484
transform 1 0 23000 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_250
timestamp 1666464484
transform 1 0 24104 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_254
timestamp 1666464484
transform 1 0 24472 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_256
timestamp 1666464484
transform 1 0 24656 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_268
timestamp 1666464484
transform 1 0 25760 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_280
timestamp 1666464484
transform 1 0 26864 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_284
timestamp 1666464484
transform 1 0 27232 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_286
timestamp 1666464484
transform 1 0 27416 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_298
timestamp 1666464484
transform 1 0 28520 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_310
timestamp 1666464484
transform 1 0 29624 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_314
timestamp 1666464484
transform 1 0 29992 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_316
timestamp 1666464484
transform 1 0 30176 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_328
timestamp 1666464484
transform 1 0 31280 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_340
timestamp 1666464484
transform 1 0 32384 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_344
timestamp 1666464484
transform 1 0 32752 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_346
timestamp 1666464484
transform 1 0 32936 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_358
timestamp 1666464484
transform 1 0 34040 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_370
timestamp 1666464484
transform 1 0 35144 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_374
timestamp 1666464484
transform 1 0 35512 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_376
timestamp 1666464484
transform 1 0 35696 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_388
timestamp 1666464484
transform 1 0 36800 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_400
timestamp 1666464484
transform 1 0 37904 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_404
timestamp 1666464484
transform 1 0 38272 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_406
timestamp 1666464484
transform 1 0 38456 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_418
timestamp 1666464484
transform 1 0 39560 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_430
timestamp 1666464484
transform 1 0 40664 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_434
timestamp 1666464484
transform 1 0 41032 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_436
timestamp 1666464484
transform 1 0 41216 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_448
timestamp 1666464484
transform 1 0 42320 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_460
timestamp 1666464484
transform 1 0 43424 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_464
timestamp 1666464484
transform 1 0 43792 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_466
timestamp 1666464484
transform 1 0 43976 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_478
timestamp 1666464484
transform 1 0 45080 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_490
timestamp 1666464484
transform 1 0 46184 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_494
timestamp 1666464484
transform 1 0 46552 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_496
timestamp 1666464484
transform 1 0 46736 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_508
timestamp 1666464484
transform 1 0 47840 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_520
timestamp 1666464484
transform 1 0 48944 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_524
timestamp 1666464484
transform 1 0 49312 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_526
timestamp 1666464484
transform 1 0 49496 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_538
timestamp 1666464484
transform 1 0 50600 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_550
timestamp 1666464484
transform 1 0 51704 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_554
timestamp 1666464484
transform 1 0 52072 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_556
timestamp 1666464484
transform 1 0 52256 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_568
timestamp 1666464484
transform 1 0 53360 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_580
timestamp 1666464484
transform 1 0 54464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_584
timestamp 1666464484
transform 1 0 54832 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_586
timestamp 1666464484
transform 1 0 55016 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_598
timestamp 1666464484
transform 1 0 56120 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_610
timestamp 1666464484
transform 1 0 57224 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_614
timestamp 1666464484
transform 1 0 57592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_616
timestamp 1666464484
transform 1 0 57776 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_624
timestamp 1666464484
transform 1 0 58512 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1666464484
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1666464484
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_27
timestamp 1666464484
transform 1 0 3588 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_31
timestamp 1666464484
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_43
timestamp 1666464484
transform 1 0 5060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_55
timestamp 1666464484
transform 1 0 6164 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_59
timestamp 1666464484
transform 1 0 6532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_61
timestamp 1666464484
transform 1 0 6716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_73
timestamp 1666464484
transform 1 0 7820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_85
timestamp 1666464484
transform 1 0 8924 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_89
timestamp 1666464484
transform 1 0 9292 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_91
timestamp 1666464484
transform 1 0 9476 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_103
timestamp 1666464484
transform 1 0 10580 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_115
timestamp 1666464484
transform 1 0 11684 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_119
timestamp 1666464484
transform 1 0 12052 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_121
timestamp 1666464484
transform 1 0 12236 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_133
timestamp 1666464484
transform 1 0 13340 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_145
timestamp 1666464484
transform 1 0 14444 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_149
timestamp 1666464484
transform 1 0 14812 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_151
timestamp 1666464484
transform 1 0 14996 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_163
timestamp 1666464484
transform 1 0 16100 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_175
timestamp 1666464484
transform 1 0 17204 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_179
timestamp 1666464484
transform 1 0 17572 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1666464484
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1666464484
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_205
timestamp 1666464484
transform 1 0 19964 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_209
timestamp 1666464484
transform 1 0 20332 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_211
timestamp 1666464484
transform 1 0 20516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_223
timestamp 1666464484
transform 1 0 21620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_235
timestamp 1666464484
transform 1 0 22724 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_239
timestamp 1666464484
transform 1 0 23092 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_241
timestamp 1666464484
transform 1 0 23276 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_253
timestamp 1666464484
transform 1 0 24380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_265
timestamp 1666464484
transform 1 0 25484 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_269
timestamp 1666464484
transform 1 0 25852 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_271
timestamp 1666464484
transform 1 0 26036 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_283
timestamp 1666464484
transform 1 0 27140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_295
timestamp 1666464484
transform 1 0 28244 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_299
timestamp 1666464484
transform 1 0 28612 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_301
timestamp 1666464484
transform 1 0 28796 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_313
timestamp 1666464484
transform 1 0 29900 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_325
timestamp 1666464484
transform 1 0 31004 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_329
timestamp 1666464484
transform 1 0 31372 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_331
timestamp 1666464484
transform 1 0 31556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_343
timestamp 1666464484
transform 1 0 32660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_355
timestamp 1666464484
transform 1 0 33764 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_359
timestamp 1666464484
transform 1 0 34132 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1666464484
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1666464484
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_385
timestamp 1666464484
transform 1 0 36524 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_389
timestamp 1666464484
transform 1 0 36892 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_391
timestamp 1666464484
transform 1 0 37076 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_403
timestamp 1666464484
transform 1 0 38180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_415
timestamp 1666464484
transform 1 0 39284 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_419
timestamp 1666464484
transform 1 0 39652 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_421
timestamp 1666464484
transform 1 0 39836 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_433
timestamp 1666464484
transform 1 0 40940 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_445
timestamp 1666464484
transform 1 0 42044 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_449
timestamp 1666464484
transform 1 0 42412 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_451
timestamp 1666464484
transform 1 0 42596 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_463
timestamp 1666464484
transform 1 0 43700 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_475
timestamp 1666464484
transform 1 0 44804 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_479
timestamp 1666464484
transform 1 0 45172 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_481
timestamp 1666464484
transform 1 0 45356 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_493
timestamp 1666464484
transform 1 0 46460 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_505
timestamp 1666464484
transform 1 0 47564 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_509
timestamp 1666464484
transform 1 0 47932 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_511
timestamp 1666464484
transform 1 0 48116 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_523
timestamp 1666464484
transform 1 0 49220 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_535
timestamp 1666464484
transform 1 0 50324 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_539
timestamp 1666464484
transform 1 0 50692 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1666464484
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_553
timestamp 1666464484
transform 1 0 51980 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_565
timestamp 1666464484
transform 1 0 53084 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_569
timestamp 1666464484
transform 1 0 53452 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_571
timestamp 1666464484
transform 1 0 53636 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_583
timestamp 1666464484
transform 1 0 54740 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_595
timestamp 1666464484
transform 1 0 55844 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_599
timestamp 1666464484
transform 1 0 56212 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_601
timestamp 1666464484
transform 1 0 56396 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_613
timestamp 1666464484
transform 1 0 57500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1666464484
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_16
timestamp 1666464484
transform 1 0 2576 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_28
timestamp 1666464484
transform 1 0 3680 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_40
timestamp 1666464484
transform 1 0 4784 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_44
timestamp 1666464484
transform 1 0 5152 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_46
timestamp 1666464484
transform 1 0 5336 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_58
timestamp 1666464484
transform 1 0 6440 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_70
timestamp 1666464484
transform 1 0 7544 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_74
timestamp 1666464484
transform 1 0 7912 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_76
timestamp 1666464484
transform 1 0 8096 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_88
timestamp 1666464484
transform 1 0 9200 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_100
timestamp 1666464484
transform 1 0 10304 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_104
timestamp 1666464484
transform 1 0 10672 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_106
timestamp 1666464484
transform 1 0 10856 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_118
timestamp 1666464484
transform 1 0 11960 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_130
timestamp 1666464484
transform 1 0 13064 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_134
timestamp 1666464484
transform 1 0 13432 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_136
timestamp 1666464484
transform 1 0 13616 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_148
timestamp 1666464484
transform 1 0 14720 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_160
timestamp 1666464484
transform 1 0 15824 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_164
timestamp 1666464484
transform 1 0 16192 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_166
timestamp 1666464484
transform 1 0 16376 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_178
timestamp 1666464484
transform 1 0 17480 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_190
timestamp 1666464484
transform 1 0 18584 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_194
timestamp 1666464484
transform 1 0 18952 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_196
timestamp 1666464484
transform 1 0 19136 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_208
timestamp 1666464484
transform 1 0 20240 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_220
timestamp 1666464484
transform 1 0 21344 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_224
timestamp 1666464484
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_226
timestamp 1666464484
transform 1 0 21896 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_238
timestamp 1666464484
transform 1 0 23000 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_250
timestamp 1666464484
transform 1 0 24104 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_254
timestamp 1666464484
transform 1 0 24472 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_256
timestamp 1666464484
transform 1 0 24656 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_268
timestamp 1666464484
transform 1 0 25760 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_280
timestamp 1666464484
transform 1 0 26864 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_284
timestamp 1666464484
transform 1 0 27232 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_286
timestamp 1666464484
transform 1 0 27416 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_298
timestamp 1666464484
transform 1 0 28520 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_310
timestamp 1666464484
transform 1 0 29624 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_314
timestamp 1666464484
transform 1 0 29992 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_316
timestamp 1666464484
transform 1 0 30176 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_328
timestamp 1666464484
transform 1 0 31280 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_340
timestamp 1666464484
transform 1 0 32384 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_344
timestamp 1666464484
transform 1 0 32752 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_346
timestamp 1666464484
transform 1 0 32936 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_358
timestamp 1666464484
transform 1 0 34040 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_370
timestamp 1666464484
transform 1 0 35144 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_374
timestamp 1666464484
transform 1 0 35512 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_376
timestamp 1666464484
transform 1 0 35696 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_388
timestamp 1666464484
transform 1 0 36800 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_400
timestamp 1666464484
transform 1 0 37904 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_404
timestamp 1666464484
transform 1 0 38272 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_406
timestamp 1666464484
transform 1 0 38456 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_418
timestamp 1666464484
transform 1 0 39560 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_430
timestamp 1666464484
transform 1 0 40664 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_434
timestamp 1666464484
transform 1 0 41032 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_436
timestamp 1666464484
transform 1 0 41216 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_448
timestamp 1666464484
transform 1 0 42320 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_460
timestamp 1666464484
transform 1 0 43424 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_464
timestamp 1666464484
transform 1 0 43792 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_466
timestamp 1666464484
transform 1 0 43976 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_478
timestamp 1666464484
transform 1 0 45080 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_490
timestamp 1666464484
transform 1 0 46184 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_494
timestamp 1666464484
transform 1 0 46552 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_496
timestamp 1666464484
transform 1 0 46736 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_508
timestamp 1666464484
transform 1 0 47840 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_520
timestamp 1666464484
transform 1 0 48944 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_524
timestamp 1666464484
transform 1 0 49312 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_526
timestamp 1666464484
transform 1 0 49496 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_538
timestamp 1666464484
transform 1 0 50600 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_550
timestamp 1666464484
transform 1 0 51704 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_554
timestamp 1666464484
transform 1 0 52072 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_556
timestamp 1666464484
transform 1 0 52256 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_568
timestamp 1666464484
transform 1 0 53360 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_580
timestamp 1666464484
transform 1 0 54464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_584
timestamp 1666464484
transform 1 0 54832 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_586
timestamp 1666464484
transform 1 0 55016 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_598
timestamp 1666464484
transform 1 0 56120 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_610
timestamp 1666464484
transform 1 0 57224 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_614
timestamp 1666464484
transform 1 0 57592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_616
timestamp 1666464484
transform 1 0 57776 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_624
timestamp 1666464484
transform 1 0 58512 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1666464484
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1666464484
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_27
timestamp 1666464484
transform 1 0 3588 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_31
timestamp 1666464484
transform 1 0 3956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_43
timestamp 1666464484
transform 1 0 5060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_55
timestamp 1666464484
transform 1 0 6164 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_59
timestamp 1666464484
transform 1 0 6532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_61
timestamp 1666464484
transform 1 0 6716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_73
timestamp 1666464484
transform 1 0 7820 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_85
timestamp 1666464484
transform 1 0 8924 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_89
timestamp 1666464484
transform 1 0 9292 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_91
timestamp 1666464484
transform 1 0 9476 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_103
timestamp 1666464484
transform 1 0 10580 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_115
timestamp 1666464484
transform 1 0 11684 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_119
timestamp 1666464484
transform 1 0 12052 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_121
timestamp 1666464484
transform 1 0 12236 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_133
timestamp 1666464484
transform 1 0 13340 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_145
timestamp 1666464484
transform 1 0 14444 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_149
timestamp 1666464484
transform 1 0 14812 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_151
timestamp 1666464484
transform 1 0 14996 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_163
timestamp 1666464484
transform 1 0 16100 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_175
timestamp 1666464484
transform 1 0 17204 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_179
timestamp 1666464484
transform 1 0 17572 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1666464484
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1666464484
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_205
timestamp 1666464484
transform 1 0 19964 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_209
timestamp 1666464484
transform 1 0 20332 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_211
timestamp 1666464484
transform 1 0 20516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_223
timestamp 1666464484
transform 1 0 21620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_235
timestamp 1666464484
transform 1 0 22724 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_239
timestamp 1666464484
transform 1 0 23092 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_241
timestamp 1666464484
transform 1 0 23276 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_253
timestamp 1666464484
transform 1 0 24380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_265
timestamp 1666464484
transform 1 0 25484 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_269
timestamp 1666464484
transform 1 0 25852 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_271
timestamp 1666464484
transform 1 0 26036 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_283
timestamp 1666464484
transform 1 0 27140 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_295
timestamp 1666464484
transform 1 0 28244 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_299
timestamp 1666464484
transform 1 0 28612 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_301
timestamp 1666464484
transform 1 0 28796 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_313
timestamp 1666464484
transform 1 0 29900 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_325
timestamp 1666464484
transform 1 0 31004 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_329
timestamp 1666464484
transform 1 0 31372 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_331
timestamp 1666464484
transform 1 0 31556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_343
timestamp 1666464484
transform 1 0 32660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_355
timestamp 1666464484
transform 1 0 33764 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_359
timestamp 1666464484
transform 1 0 34132 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1666464484
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1666464484
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_385
timestamp 1666464484
transform 1 0 36524 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_389
timestamp 1666464484
transform 1 0 36892 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_391
timestamp 1666464484
transform 1 0 37076 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_403
timestamp 1666464484
transform 1 0 38180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_415
timestamp 1666464484
transform 1 0 39284 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_419
timestamp 1666464484
transform 1 0 39652 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_421
timestamp 1666464484
transform 1 0 39836 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_433
timestamp 1666464484
transform 1 0 40940 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_445
timestamp 1666464484
transform 1 0 42044 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_449
timestamp 1666464484
transform 1 0 42412 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_451
timestamp 1666464484
transform 1 0 42596 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_463
timestamp 1666464484
transform 1 0 43700 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_475
timestamp 1666464484
transform 1 0 44804 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_479
timestamp 1666464484
transform 1 0 45172 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_481
timestamp 1666464484
transform 1 0 45356 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_493
timestamp 1666464484
transform 1 0 46460 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_505
timestamp 1666464484
transform 1 0 47564 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_509
timestamp 1666464484
transform 1 0 47932 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_511
timestamp 1666464484
transform 1 0 48116 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_523
timestamp 1666464484
transform 1 0 49220 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_535
timestamp 1666464484
transform 1 0 50324 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_539
timestamp 1666464484
transform 1 0 50692 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1666464484
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_553
timestamp 1666464484
transform 1 0 51980 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_565
timestamp 1666464484
transform 1 0 53084 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_569
timestamp 1666464484
transform 1 0 53452 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_571
timestamp 1666464484
transform 1 0 53636 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_583
timestamp 1666464484
transform 1 0 54740 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_595
timestamp 1666464484
transform 1 0 55844 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_599
timestamp 1666464484
transform 1 0 56212 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_601
timestamp 1666464484
transform 1 0 56396 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_613
timestamp 1666464484
transform 1 0 57500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1666464484
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_16
timestamp 1666464484
transform 1 0 2576 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_28
timestamp 1666464484
transform 1 0 3680 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_40
timestamp 1666464484
transform 1 0 4784 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_44
timestamp 1666464484
transform 1 0 5152 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_46
timestamp 1666464484
transform 1 0 5336 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_58
timestamp 1666464484
transform 1 0 6440 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_70
timestamp 1666464484
transform 1 0 7544 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_74
timestamp 1666464484
transform 1 0 7912 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_76
timestamp 1666464484
transform 1 0 8096 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_88
timestamp 1666464484
transform 1 0 9200 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_100
timestamp 1666464484
transform 1 0 10304 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_104
timestamp 1666464484
transform 1 0 10672 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_106
timestamp 1666464484
transform 1 0 10856 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_118
timestamp 1666464484
transform 1 0 11960 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_130
timestamp 1666464484
transform 1 0 13064 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_134
timestamp 1666464484
transform 1 0 13432 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_136
timestamp 1666464484
transform 1 0 13616 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_148
timestamp 1666464484
transform 1 0 14720 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_160
timestamp 1666464484
transform 1 0 15824 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_164
timestamp 1666464484
transform 1 0 16192 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_166
timestamp 1666464484
transform 1 0 16376 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_178
timestamp 1666464484
transform 1 0 17480 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_190
timestamp 1666464484
transform 1 0 18584 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_194
timestamp 1666464484
transform 1 0 18952 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_196
timestamp 1666464484
transform 1 0 19136 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_208
timestamp 1666464484
transform 1 0 20240 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_220
timestamp 1666464484
transform 1 0 21344 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_224
timestamp 1666464484
transform 1 0 21712 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_226
timestamp 1666464484
transform 1 0 21896 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_238
timestamp 1666464484
transform 1 0 23000 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_250
timestamp 1666464484
transform 1 0 24104 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_254
timestamp 1666464484
transform 1 0 24472 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_256
timestamp 1666464484
transform 1 0 24656 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_268
timestamp 1666464484
transform 1 0 25760 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_280
timestamp 1666464484
transform 1 0 26864 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_284
timestamp 1666464484
transform 1 0 27232 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_286
timestamp 1666464484
transform 1 0 27416 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_298
timestamp 1666464484
transform 1 0 28520 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_310
timestamp 1666464484
transform 1 0 29624 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_314
timestamp 1666464484
transform 1 0 29992 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_316
timestamp 1666464484
transform 1 0 30176 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_328
timestamp 1666464484
transform 1 0 31280 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_340
timestamp 1666464484
transform 1 0 32384 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_344
timestamp 1666464484
transform 1 0 32752 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_346
timestamp 1666464484
transform 1 0 32936 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_358
timestamp 1666464484
transform 1 0 34040 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_370
timestamp 1666464484
transform 1 0 35144 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_374
timestamp 1666464484
transform 1 0 35512 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_376
timestamp 1666464484
transform 1 0 35696 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_388
timestamp 1666464484
transform 1 0 36800 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_400
timestamp 1666464484
transform 1 0 37904 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_404
timestamp 1666464484
transform 1 0 38272 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_406
timestamp 1666464484
transform 1 0 38456 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_418
timestamp 1666464484
transform 1 0 39560 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_430
timestamp 1666464484
transform 1 0 40664 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_434
timestamp 1666464484
transform 1 0 41032 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_436
timestamp 1666464484
transform 1 0 41216 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_448
timestamp 1666464484
transform 1 0 42320 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_460
timestamp 1666464484
transform 1 0 43424 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_464
timestamp 1666464484
transform 1 0 43792 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_466
timestamp 1666464484
transform 1 0 43976 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_478
timestamp 1666464484
transform 1 0 45080 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_490
timestamp 1666464484
transform 1 0 46184 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_494
timestamp 1666464484
transform 1 0 46552 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_496
timestamp 1666464484
transform 1 0 46736 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_508
timestamp 1666464484
transform 1 0 47840 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_520
timestamp 1666464484
transform 1 0 48944 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_524
timestamp 1666464484
transform 1 0 49312 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_526
timestamp 1666464484
transform 1 0 49496 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_538
timestamp 1666464484
transform 1 0 50600 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_550
timestamp 1666464484
transform 1 0 51704 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_554
timestamp 1666464484
transform 1 0 52072 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_556
timestamp 1666464484
transform 1 0 52256 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_568
timestamp 1666464484
transform 1 0 53360 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_580
timestamp 1666464484
transform 1 0 54464 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_584
timestamp 1666464484
transform 1 0 54832 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_586
timestamp 1666464484
transform 1 0 55016 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_598
timestamp 1666464484
transform 1 0 56120 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_610
timestamp 1666464484
transform 1 0 57224 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_614
timestamp 1666464484
transform 1 0 57592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_616
timestamp 1666464484
transform 1 0 57776 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_624
timestamp 1666464484
transform 1 0 58512 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1666464484
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1666464484
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_27
timestamp 1666464484
transform 1 0 3588 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_31
timestamp 1666464484
transform 1 0 3956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_43
timestamp 1666464484
transform 1 0 5060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_55
timestamp 1666464484
transform 1 0 6164 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_59
timestamp 1666464484
transform 1 0 6532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_61
timestamp 1666464484
transform 1 0 6716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_73
timestamp 1666464484
transform 1 0 7820 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_85
timestamp 1666464484
transform 1 0 8924 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_89
timestamp 1666464484
transform 1 0 9292 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_91
timestamp 1666464484
transform 1 0 9476 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_103
timestamp 1666464484
transform 1 0 10580 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_115
timestamp 1666464484
transform 1 0 11684 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_119
timestamp 1666464484
transform 1 0 12052 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_121
timestamp 1666464484
transform 1 0 12236 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_133
timestamp 1666464484
transform 1 0 13340 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_145
timestamp 1666464484
transform 1 0 14444 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_149
timestamp 1666464484
transform 1 0 14812 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_151
timestamp 1666464484
transform 1 0 14996 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_163
timestamp 1666464484
transform 1 0 16100 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_175
timestamp 1666464484
transform 1 0 17204 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_179
timestamp 1666464484
transform 1 0 17572 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1666464484
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1666464484
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_205
timestamp 1666464484
transform 1 0 19964 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_209
timestamp 1666464484
transform 1 0 20332 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_211
timestamp 1666464484
transform 1 0 20516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_223
timestamp 1666464484
transform 1 0 21620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_235
timestamp 1666464484
transform 1 0 22724 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_239
timestamp 1666464484
transform 1 0 23092 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_241
timestamp 1666464484
transform 1 0 23276 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_253
timestamp 1666464484
transform 1 0 24380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_265
timestamp 1666464484
transform 1 0 25484 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_269
timestamp 1666464484
transform 1 0 25852 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_271
timestamp 1666464484
transform 1 0 26036 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_283
timestamp 1666464484
transform 1 0 27140 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_295
timestamp 1666464484
transform 1 0 28244 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_299
timestamp 1666464484
transform 1 0 28612 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_301
timestamp 1666464484
transform 1 0 28796 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_313
timestamp 1666464484
transform 1 0 29900 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_325
timestamp 1666464484
transform 1 0 31004 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_329
timestamp 1666464484
transform 1 0 31372 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_331
timestamp 1666464484
transform 1 0 31556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_343
timestamp 1666464484
transform 1 0 32660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_355
timestamp 1666464484
transform 1 0 33764 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_359
timestamp 1666464484
transform 1 0 34132 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1666464484
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1666464484
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_385
timestamp 1666464484
transform 1 0 36524 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_389
timestamp 1666464484
transform 1 0 36892 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_391
timestamp 1666464484
transform 1 0 37076 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_403
timestamp 1666464484
transform 1 0 38180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_415
timestamp 1666464484
transform 1 0 39284 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_419
timestamp 1666464484
transform 1 0 39652 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_421
timestamp 1666464484
transform 1 0 39836 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_433
timestamp 1666464484
transform 1 0 40940 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_445
timestamp 1666464484
transform 1 0 42044 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_449
timestamp 1666464484
transform 1 0 42412 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_451
timestamp 1666464484
transform 1 0 42596 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_463
timestamp 1666464484
transform 1 0 43700 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_475
timestamp 1666464484
transform 1 0 44804 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_479
timestamp 1666464484
transform 1 0 45172 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_481
timestamp 1666464484
transform 1 0 45356 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_493
timestamp 1666464484
transform 1 0 46460 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_505
timestamp 1666464484
transform 1 0 47564 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_509
timestamp 1666464484
transform 1 0 47932 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_511
timestamp 1666464484
transform 1 0 48116 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_523
timestamp 1666464484
transform 1 0 49220 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_535
timestamp 1666464484
transform 1 0 50324 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_539
timestamp 1666464484
transform 1 0 50692 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1666464484
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_553
timestamp 1666464484
transform 1 0 51980 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_565
timestamp 1666464484
transform 1 0 53084 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_569
timestamp 1666464484
transform 1 0 53452 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_571
timestamp 1666464484
transform 1 0 53636 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_583
timestamp 1666464484
transform 1 0 54740 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_595
timestamp 1666464484
transform 1 0 55844 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_599
timestamp 1666464484
transform 1 0 56212 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_601
timestamp 1666464484
transform 1 0 56396 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_613
timestamp 1666464484
transform 1 0 57500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1666464484
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_16
timestamp 1666464484
transform 1 0 2576 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_28
timestamp 1666464484
transform 1 0 3680 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_40
timestamp 1666464484
transform 1 0 4784 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_44
timestamp 1666464484
transform 1 0 5152 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_46
timestamp 1666464484
transform 1 0 5336 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_58
timestamp 1666464484
transform 1 0 6440 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_70
timestamp 1666464484
transform 1 0 7544 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_74
timestamp 1666464484
transform 1 0 7912 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_76
timestamp 1666464484
transform 1 0 8096 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_88
timestamp 1666464484
transform 1 0 9200 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_100
timestamp 1666464484
transform 1 0 10304 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_104
timestamp 1666464484
transform 1 0 10672 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_106
timestamp 1666464484
transform 1 0 10856 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_118
timestamp 1666464484
transform 1 0 11960 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_130
timestamp 1666464484
transform 1 0 13064 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_134
timestamp 1666464484
transform 1 0 13432 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_136
timestamp 1666464484
transform 1 0 13616 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_148
timestamp 1666464484
transform 1 0 14720 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_160
timestamp 1666464484
transform 1 0 15824 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_164
timestamp 1666464484
transform 1 0 16192 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_166
timestamp 1666464484
transform 1 0 16376 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_178
timestamp 1666464484
transform 1 0 17480 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_190
timestamp 1666464484
transform 1 0 18584 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_194
timestamp 1666464484
transform 1 0 18952 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_196
timestamp 1666464484
transform 1 0 19136 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_208
timestamp 1666464484
transform 1 0 20240 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_220
timestamp 1666464484
transform 1 0 21344 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_224
timestamp 1666464484
transform 1 0 21712 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_226
timestamp 1666464484
transform 1 0 21896 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_238
timestamp 1666464484
transform 1 0 23000 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_250
timestamp 1666464484
transform 1 0 24104 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_254
timestamp 1666464484
transform 1 0 24472 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_256
timestamp 1666464484
transform 1 0 24656 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_268
timestamp 1666464484
transform 1 0 25760 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_280
timestamp 1666464484
transform 1 0 26864 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_284
timestamp 1666464484
transform 1 0 27232 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_286
timestamp 1666464484
transform 1 0 27416 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_298
timestamp 1666464484
transform 1 0 28520 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_310
timestamp 1666464484
transform 1 0 29624 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_314
timestamp 1666464484
transform 1 0 29992 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_316
timestamp 1666464484
transform 1 0 30176 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_328
timestamp 1666464484
transform 1 0 31280 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_340
timestamp 1666464484
transform 1 0 32384 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_344
timestamp 1666464484
transform 1 0 32752 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_346
timestamp 1666464484
transform 1 0 32936 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_358
timestamp 1666464484
transform 1 0 34040 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_370
timestamp 1666464484
transform 1 0 35144 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_374
timestamp 1666464484
transform 1 0 35512 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_376
timestamp 1666464484
transform 1 0 35696 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_388
timestamp 1666464484
transform 1 0 36800 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_400
timestamp 1666464484
transform 1 0 37904 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_404
timestamp 1666464484
transform 1 0 38272 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_406
timestamp 1666464484
transform 1 0 38456 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_418
timestamp 1666464484
transform 1 0 39560 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_430
timestamp 1666464484
transform 1 0 40664 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_434
timestamp 1666464484
transform 1 0 41032 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_436
timestamp 1666464484
transform 1 0 41216 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_448
timestamp 1666464484
transform 1 0 42320 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_460
timestamp 1666464484
transform 1 0 43424 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_464
timestamp 1666464484
transform 1 0 43792 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_466
timestamp 1666464484
transform 1 0 43976 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_478
timestamp 1666464484
transform 1 0 45080 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_490
timestamp 1666464484
transform 1 0 46184 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_494
timestamp 1666464484
transform 1 0 46552 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_496
timestamp 1666464484
transform 1 0 46736 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_508
timestamp 1666464484
transform 1 0 47840 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_520
timestamp 1666464484
transform 1 0 48944 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_524
timestamp 1666464484
transform 1 0 49312 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_526
timestamp 1666464484
transform 1 0 49496 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_538
timestamp 1666464484
transform 1 0 50600 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_550
timestamp 1666464484
transform 1 0 51704 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_554
timestamp 1666464484
transform 1 0 52072 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_556
timestamp 1666464484
transform 1 0 52256 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_568
timestamp 1666464484
transform 1 0 53360 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_580
timestamp 1666464484
transform 1 0 54464 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_584
timestamp 1666464484
transform 1 0 54832 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_586
timestamp 1666464484
transform 1 0 55016 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_598
timestamp 1666464484
transform 1 0 56120 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_610
timestamp 1666464484
transform 1 0 57224 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_614
timestamp 1666464484
transform 1 0 57592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_616
timestamp 1666464484
transform 1 0 57776 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_624
timestamp 1666464484
transform 1 0 58512 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1666464484
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1666464484
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_27
timestamp 1666464484
transform 1 0 3588 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_31
timestamp 1666464484
transform 1 0 3956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_43
timestamp 1666464484
transform 1 0 5060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_55
timestamp 1666464484
transform 1 0 6164 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_59
timestamp 1666464484
transform 1 0 6532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_61
timestamp 1666464484
transform 1 0 6716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_73
timestamp 1666464484
transform 1 0 7820 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_85
timestamp 1666464484
transform 1 0 8924 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_89
timestamp 1666464484
transform 1 0 9292 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_91
timestamp 1666464484
transform 1 0 9476 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_103
timestamp 1666464484
transform 1 0 10580 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_115
timestamp 1666464484
transform 1 0 11684 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_119
timestamp 1666464484
transform 1 0 12052 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_121
timestamp 1666464484
transform 1 0 12236 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_133
timestamp 1666464484
transform 1 0 13340 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_145
timestamp 1666464484
transform 1 0 14444 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_149
timestamp 1666464484
transform 1 0 14812 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_151
timestamp 1666464484
transform 1 0 14996 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_163
timestamp 1666464484
transform 1 0 16100 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_175
timestamp 1666464484
transform 1 0 17204 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_179
timestamp 1666464484
transform 1 0 17572 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1666464484
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1666464484
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_205
timestamp 1666464484
transform 1 0 19964 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_209
timestamp 1666464484
transform 1 0 20332 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_211
timestamp 1666464484
transform 1 0 20516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_223
timestamp 1666464484
transform 1 0 21620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_235
timestamp 1666464484
transform 1 0 22724 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_239
timestamp 1666464484
transform 1 0 23092 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_241
timestamp 1666464484
transform 1 0 23276 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_253
timestamp 1666464484
transform 1 0 24380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_265
timestamp 1666464484
transform 1 0 25484 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_269
timestamp 1666464484
transform 1 0 25852 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_271
timestamp 1666464484
transform 1 0 26036 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_283
timestamp 1666464484
transform 1 0 27140 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_295
timestamp 1666464484
transform 1 0 28244 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_299
timestamp 1666464484
transform 1 0 28612 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_301
timestamp 1666464484
transform 1 0 28796 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_313
timestamp 1666464484
transform 1 0 29900 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_325
timestamp 1666464484
transform 1 0 31004 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_329
timestamp 1666464484
transform 1 0 31372 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_331
timestamp 1666464484
transform 1 0 31556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_343
timestamp 1666464484
transform 1 0 32660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_355
timestamp 1666464484
transform 1 0 33764 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_359
timestamp 1666464484
transform 1 0 34132 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1666464484
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1666464484
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_385
timestamp 1666464484
transform 1 0 36524 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_389
timestamp 1666464484
transform 1 0 36892 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_391
timestamp 1666464484
transform 1 0 37076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_403
timestamp 1666464484
transform 1 0 38180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_415
timestamp 1666464484
transform 1 0 39284 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_419
timestamp 1666464484
transform 1 0 39652 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_421
timestamp 1666464484
transform 1 0 39836 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_433
timestamp 1666464484
transform 1 0 40940 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_445
timestamp 1666464484
transform 1 0 42044 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_449
timestamp 1666464484
transform 1 0 42412 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_451
timestamp 1666464484
transform 1 0 42596 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_463
timestamp 1666464484
transform 1 0 43700 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_475
timestamp 1666464484
transform 1 0 44804 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_479
timestamp 1666464484
transform 1 0 45172 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_481
timestamp 1666464484
transform 1 0 45356 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_493
timestamp 1666464484
transform 1 0 46460 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_505
timestamp 1666464484
transform 1 0 47564 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_509
timestamp 1666464484
transform 1 0 47932 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_511
timestamp 1666464484
transform 1 0 48116 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_523
timestamp 1666464484
transform 1 0 49220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_535
timestamp 1666464484
transform 1 0 50324 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_539
timestamp 1666464484
transform 1 0 50692 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1666464484
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_553
timestamp 1666464484
transform 1 0 51980 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_565
timestamp 1666464484
transform 1 0 53084 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_569
timestamp 1666464484
transform 1 0 53452 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_571
timestamp 1666464484
transform 1 0 53636 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_583
timestamp 1666464484
transform 1 0 54740 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_595
timestamp 1666464484
transform 1 0 55844 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_599
timestamp 1666464484
transform 1 0 56212 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_601
timestamp 1666464484
transform 1 0 56396 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_613
timestamp 1666464484
transform 1 0 57500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1666464484
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_16
timestamp 1666464484
transform 1 0 2576 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_28
timestamp 1666464484
transform 1 0 3680 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_40
timestamp 1666464484
transform 1 0 4784 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_44
timestamp 1666464484
transform 1 0 5152 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_46
timestamp 1666464484
transform 1 0 5336 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_58
timestamp 1666464484
transform 1 0 6440 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_70
timestamp 1666464484
transform 1 0 7544 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_74
timestamp 1666464484
transform 1 0 7912 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_76
timestamp 1666464484
transform 1 0 8096 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_88
timestamp 1666464484
transform 1 0 9200 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_100
timestamp 1666464484
transform 1 0 10304 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_104
timestamp 1666464484
transform 1 0 10672 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_106
timestamp 1666464484
transform 1 0 10856 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_118
timestamp 1666464484
transform 1 0 11960 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_130
timestamp 1666464484
transform 1 0 13064 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_134
timestamp 1666464484
transform 1 0 13432 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_136
timestamp 1666464484
transform 1 0 13616 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_148
timestamp 1666464484
transform 1 0 14720 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_160
timestamp 1666464484
transform 1 0 15824 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_164
timestamp 1666464484
transform 1 0 16192 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_166
timestamp 1666464484
transform 1 0 16376 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_178
timestamp 1666464484
transform 1 0 17480 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_190
timestamp 1666464484
transform 1 0 18584 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_194
timestamp 1666464484
transform 1 0 18952 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_196
timestamp 1666464484
transform 1 0 19136 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_208
timestamp 1666464484
transform 1 0 20240 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_220
timestamp 1666464484
transform 1 0 21344 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_224
timestamp 1666464484
transform 1 0 21712 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_226
timestamp 1666464484
transform 1 0 21896 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_238
timestamp 1666464484
transform 1 0 23000 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_250
timestamp 1666464484
transform 1 0 24104 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_254
timestamp 1666464484
transform 1 0 24472 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_256
timestamp 1666464484
transform 1 0 24656 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_268
timestamp 1666464484
transform 1 0 25760 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_280
timestamp 1666464484
transform 1 0 26864 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_284
timestamp 1666464484
transform 1 0 27232 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_286
timestamp 1666464484
transform 1 0 27416 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_298
timestamp 1666464484
transform 1 0 28520 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_310
timestamp 1666464484
transform 1 0 29624 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_314
timestamp 1666464484
transform 1 0 29992 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_316
timestamp 1666464484
transform 1 0 30176 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_328
timestamp 1666464484
transform 1 0 31280 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_340
timestamp 1666464484
transform 1 0 32384 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_344
timestamp 1666464484
transform 1 0 32752 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_346
timestamp 1666464484
transform 1 0 32936 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_358
timestamp 1666464484
transform 1 0 34040 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_370
timestamp 1666464484
transform 1 0 35144 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_374
timestamp 1666464484
transform 1 0 35512 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_376
timestamp 1666464484
transform 1 0 35696 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_388
timestamp 1666464484
transform 1 0 36800 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_400
timestamp 1666464484
transform 1 0 37904 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_404
timestamp 1666464484
transform 1 0 38272 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_406
timestamp 1666464484
transform 1 0 38456 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_418
timestamp 1666464484
transform 1 0 39560 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_430
timestamp 1666464484
transform 1 0 40664 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_434
timestamp 1666464484
transform 1 0 41032 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_436
timestamp 1666464484
transform 1 0 41216 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_448
timestamp 1666464484
transform 1 0 42320 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_460
timestamp 1666464484
transform 1 0 43424 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_464
timestamp 1666464484
transform 1 0 43792 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_466
timestamp 1666464484
transform 1 0 43976 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_478
timestamp 1666464484
transform 1 0 45080 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_490
timestamp 1666464484
transform 1 0 46184 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_494
timestamp 1666464484
transform 1 0 46552 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_496
timestamp 1666464484
transform 1 0 46736 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_508
timestamp 1666464484
transform 1 0 47840 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_520
timestamp 1666464484
transform 1 0 48944 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_524
timestamp 1666464484
transform 1 0 49312 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_526
timestamp 1666464484
transform 1 0 49496 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_538
timestamp 1666464484
transform 1 0 50600 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_550
timestamp 1666464484
transform 1 0 51704 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_554
timestamp 1666464484
transform 1 0 52072 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_556
timestamp 1666464484
transform 1 0 52256 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_568
timestamp 1666464484
transform 1 0 53360 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_580
timestamp 1666464484
transform 1 0 54464 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_584
timestamp 1666464484
transform 1 0 54832 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_586
timestamp 1666464484
transform 1 0 55016 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_598
timestamp 1666464484
transform 1 0 56120 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_610
timestamp 1666464484
transform 1 0 57224 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_614
timestamp 1666464484
transform 1 0 57592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_616
timestamp 1666464484
transform 1 0 57776 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_624
timestamp 1666464484
transform 1 0 58512 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1666464484
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1666464484
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_27
timestamp 1666464484
transform 1 0 3588 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_31
timestamp 1666464484
transform 1 0 3956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_43
timestamp 1666464484
transform 1 0 5060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_55
timestamp 1666464484
transform 1 0 6164 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_59
timestamp 1666464484
transform 1 0 6532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_61
timestamp 1666464484
transform 1 0 6716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_73
timestamp 1666464484
transform 1 0 7820 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_85
timestamp 1666464484
transform 1 0 8924 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_89
timestamp 1666464484
transform 1 0 9292 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_91
timestamp 1666464484
transform 1 0 9476 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_103
timestamp 1666464484
transform 1 0 10580 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_115
timestamp 1666464484
transform 1 0 11684 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_119
timestamp 1666464484
transform 1 0 12052 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_121
timestamp 1666464484
transform 1 0 12236 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_133
timestamp 1666464484
transform 1 0 13340 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_145
timestamp 1666464484
transform 1 0 14444 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_149
timestamp 1666464484
transform 1 0 14812 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_151
timestamp 1666464484
transform 1 0 14996 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_163
timestamp 1666464484
transform 1 0 16100 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_175
timestamp 1666464484
transform 1 0 17204 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_179
timestamp 1666464484
transform 1 0 17572 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1666464484
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1666464484
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_205
timestamp 1666464484
transform 1 0 19964 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_209
timestamp 1666464484
transform 1 0 20332 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_211
timestamp 1666464484
transform 1 0 20516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_223
timestamp 1666464484
transform 1 0 21620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_235
timestamp 1666464484
transform 1 0 22724 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_239
timestamp 1666464484
transform 1 0 23092 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_241
timestamp 1666464484
transform 1 0 23276 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_253
timestamp 1666464484
transform 1 0 24380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_265
timestamp 1666464484
transform 1 0 25484 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_269
timestamp 1666464484
transform 1 0 25852 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_271
timestamp 1666464484
transform 1 0 26036 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_283
timestamp 1666464484
transform 1 0 27140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_295
timestamp 1666464484
transform 1 0 28244 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_299
timestamp 1666464484
transform 1 0 28612 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_301
timestamp 1666464484
transform 1 0 28796 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_313
timestamp 1666464484
transform 1 0 29900 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_325
timestamp 1666464484
transform 1 0 31004 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_329
timestamp 1666464484
transform 1 0 31372 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_331
timestamp 1666464484
transform 1 0 31556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_343
timestamp 1666464484
transform 1 0 32660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_355
timestamp 1666464484
transform 1 0 33764 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_359
timestamp 1666464484
transform 1 0 34132 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1666464484
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1666464484
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_385
timestamp 1666464484
transform 1 0 36524 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_389
timestamp 1666464484
transform 1 0 36892 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_391
timestamp 1666464484
transform 1 0 37076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_403
timestamp 1666464484
transform 1 0 38180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_415
timestamp 1666464484
transform 1 0 39284 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_419
timestamp 1666464484
transform 1 0 39652 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_421
timestamp 1666464484
transform 1 0 39836 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_433
timestamp 1666464484
transform 1 0 40940 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_445
timestamp 1666464484
transform 1 0 42044 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_449
timestamp 1666464484
transform 1 0 42412 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_451
timestamp 1666464484
transform 1 0 42596 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_463
timestamp 1666464484
transform 1 0 43700 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_475
timestamp 1666464484
transform 1 0 44804 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_479
timestamp 1666464484
transform 1 0 45172 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_481
timestamp 1666464484
transform 1 0 45356 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_493
timestamp 1666464484
transform 1 0 46460 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_505
timestamp 1666464484
transform 1 0 47564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_509
timestamp 1666464484
transform 1 0 47932 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_511
timestamp 1666464484
transform 1 0 48116 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_523
timestamp 1666464484
transform 1 0 49220 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_535
timestamp 1666464484
transform 1 0 50324 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_539
timestamp 1666464484
transform 1 0 50692 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1666464484
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_553
timestamp 1666464484
transform 1 0 51980 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_565
timestamp 1666464484
transform 1 0 53084 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_569
timestamp 1666464484
transform 1 0 53452 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_571
timestamp 1666464484
transform 1 0 53636 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_583
timestamp 1666464484
transform 1 0 54740 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_595
timestamp 1666464484
transform 1 0 55844 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_599
timestamp 1666464484
transform 1 0 56212 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_601
timestamp 1666464484
transform 1 0 56396 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_613
timestamp 1666464484
transform 1 0 57500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1666464484
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_16
timestamp 1666464484
transform 1 0 2576 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_28
timestamp 1666464484
transform 1 0 3680 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_40
timestamp 1666464484
transform 1 0 4784 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_44
timestamp 1666464484
transform 1 0 5152 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_46
timestamp 1666464484
transform 1 0 5336 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_58
timestamp 1666464484
transform 1 0 6440 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_70
timestamp 1666464484
transform 1 0 7544 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_74
timestamp 1666464484
transform 1 0 7912 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_76
timestamp 1666464484
transform 1 0 8096 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_88
timestamp 1666464484
transform 1 0 9200 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_100
timestamp 1666464484
transform 1 0 10304 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_104
timestamp 1666464484
transform 1 0 10672 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_106
timestamp 1666464484
transform 1 0 10856 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_118
timestamp 1666464484
transform 1 0 11960 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_130
timestamp 1666464484
transform 1 0 13064 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_134
timestamp 1666464484
transform 1 0 13432 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_136
timestamp 1666464484
transform 1 0 13616 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_148
timestamp 1666464484
transform 1 0 14720 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_160
timestamp 1666464484
transform 1 0 15824 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_164
timestamp 1666464484
transform 1 0 16192 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_166
timestamp 1666464484
transform 1 0 16376 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_178
timestamp 1666464484
transform 1 0 17480 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_190
timestamp 1666464484
transform 1 0 18584 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_194
timestamp 1666464484
transform 1 0 18952 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_196
timestamp 1666464484
transform 1 0 19136 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_208
timestamp 1666464484
transform 1 0 20240 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_220
timestamp 1666464484
transform 1 0 21344 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_224
timestamp 1666464484
transform 1 0 21712 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_226
timestamp 1666464484
transform 1 0 21896 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_238
timestamp 1666464484
transform 1 0 23000 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_250
timestamp 1666464484
transform 1 0 24104 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_254
timestamp 1666464484
transform 1 0 24472 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_256
timestamp 1666464484
transform 1 0 24656 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_268
timestamp 1666464484
transform 1 0 25760 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_280
timestamp 1666464484
transform 1 0 26864 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_284
timestamp 1666464484
transform 1 0 27232 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_286
timestamp 1666464484
transform 1 0 27416 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_298
timestamp 1666464484
transform 1 0 28520 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_310
timestamp 1666464484
transform 1 0 29624 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_314
timestamp 1666464484
transform 1 0 29992 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_316
timestamp 1666464484
transform 1 0 30176 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_328
timestamp 1666464484
transform 1 0 31280 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_340
timestamp 1666464484
transform 1 0 32384 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_344
timestamp 1666464484
transform 1 0 32752 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_346
timestamp 1666464484
transform 1 0 32936 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_358
timestamp 1666464484
transform 1 0 34040 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_370
timestamp 1666464484
transform 1 0 35144 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_374
timestamp 1666464484
transform 1 0 35512 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_376
timestamp 1666464484
transform 1 0 35696 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_388
timestamp 1666464484
transform 1 0 36800 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_400
timestamp 1666464484
transform 1 0 37904 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_404
timestamp 1666464484
transform 1 0 38272 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_406
timestamp 1666464484
transform 1 0 38456 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_418
timestamp 1666464484
transform 1 0 39560 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_430
timestamp 1666464484
transform 1 0 40664 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_434
timestamp 1666464484
transform 1 0 41032 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_436
timestamp 1666464484
transform 1 0 41216 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_448
timestamp 1666464484
transform 1 0 42320 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_460
timestamp 1666464484
transform 1 0 43424 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_464
timestamp 1666464484
transform 1 0 43792 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_466
timestamp 1666464484
transform 1 0 43976 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_478
timestamp 1666464484
transform 1 0 45080 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_490
timestamp 1666464484
transform 1 0 46184 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_494
timestamp 1666464484
transform 1 0 46552 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_496
timestamp 1666464484
transform 1 0 46736 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_508
timestamp 1666464484
transform 1 0 47840 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_520
timestamp 1666464484
transform 1 0 48944 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_524
timestamp 1666464484
transform 1 0 49312 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_526
timestamp 1666464484
transform 1 0 49496 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_538
timestamp 1666464484
transform 1 0 50600 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_550
timestamp 1666464484
transform 1 0 51704 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_554
timestamp 1666464484
transform 1 0 52072 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_556
timestamp 1666464484
transform 1 0 52256 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_568
timestamp 1666464484
transform 1 0 53360 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_580
timestamp 1666464484
transform 1 0 54464 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_584
timestamp 1666464484
transform 1 0 54832 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_586
timestamp 1666464484
transform 1 0 55016 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_598
timestamp 1666464484
transform 1 0 56120 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_610
timestamp 1666464484
transform 1 0 57224 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_614
timestamp 1666464484
transform 1 0 57592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_616
timestamp 1666464484
transform 1 0 57776 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_624
timestamp 1666464484
transform 1 0 58512 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1666464484
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1666464484
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_27
timestamp 1666464484
transform 1 0 3588 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_31
timestamp 1666464484
transform 1 0 3956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_43
timestamp 1666464484
transform 1 0 5060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_55
timestamp 1666464484
transform 1 0 6164 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_59
timestamp 1666464484
transform 1 0 6532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_61
timestamp 1666464484
transform 1 0 6716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_73
timestamp 1666464484
transform 1 0 7820 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_85
timestamp 1666464484
transform 1 0 8924 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_89
timestamp 1666464484
transform 1 0 9292 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_91
timestamp 1666464484
transform 1 0 9476 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_103
timestamp 1666464484
transform 1 0 10580 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_115
timestamp 1666464484
transform 1 0 11684 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_119
timestamp 1666464484
transform 1 0 12052 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_121
timestamp 1666464484
transform 1 0 12236 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_133
timestamp 1666464484
transform 1 0 13340 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_145
timestamp 1666464484
transform 1 0 14444 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_149
timestamp 1666464484
transform 1 0 14812 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_151
timestamp 1666464484
transform 1 0 14996 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_163
timestamp 1666464484
transform 1 0 16100 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_175
timestamp 1666464484
transform 1 0 17204 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_179
timestamp 1666464484
transform 1 0 17572 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1666464484
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1666464484
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_205
timestamp 1666464484
transform 1 0 19964 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_209
timestamp 1666464484
transform 1 0 20332 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_211
timestamp 1666464484
transform 1 0 20516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_223
timestamp 1666464484
transform 1 0 21620 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_235
timestamp 1666464484
transform 1 0 22724 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_239
timestamp 1666464484
transform 1 0 23092 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_241
timestamp 1666464484
transform 1 0 23276 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_253
timestamp 1666464484
transform 1 0 24380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_265
timestamp 1666464484
transform 1 0 25484 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_269
timestamp 1666464484
transform 1 0 25852 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_271
timestamp 1666464484
transform 1 0 26036 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_283
timestamp 1666464484
transform 1 0 27140 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_295
timestamp 1666464484
transform 1 0 28244 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_299
timestamp 1666464484
transform 1 0 28612 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_301
timestamp 1666464484
transform 1 0 28796 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_313
timestamp 1666464484
transform 1 0 29900 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_325
timestamp 1666464484
transform 1 0 31004 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_329
timestamp 1666464484
transform 1 0 31372 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_331
timestamp 1666464484
transform 1 0 31556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_343
timestamp 1666464484
transform 1 0 32660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_355
timestamp 1666464484
transform 1 0 33764 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_359
timestamp 1666464484
transform 1 0 34132 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1666464484
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1666464484
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_385
timestamp 1666464484
transform 1 0 36524 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_389
timestamp 1666464484
transform 1 0 36892 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_391
timestamp 1666464484
transform 1 0 37076 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_403
timestamp 1666464484
transform 1 0 38180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_415
timestamp 1666464484
transform 1 0 39284 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_419
timestamp 1666464484
transform 1 0 39652 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_421
timestamp 1666464484
transform 1 0 39836 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_433
timestamp 1666464484
transform 1 0 40940 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_445
timestamp 1666464484
transform 1 0 42044 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_449
timestamp 1666464484
transform 1 0 42412 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_451
timestamp 1666464484
transform 1 0 42596 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_463
timestamp 1666464484
transform 1 0 43700 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_475
timestamp 1666464484
transform 1 0 44804 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_479
timestamp 1666464484
transform 1 0 45172 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_481
timestamp 1666464484
transform 1 0 45356 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_493
timestamp 1666464484
transform 1 0 46460 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_505
timestamp 1666464484
transform 1 0 47564 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_509
timestamp 1666464484
transform 1 0 47932 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_511
timestamp 1666464484
transform 1 0 48116 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_523
timestamp 1666464484
transform 1 0 49220 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_535
timestamp 1666464484
transform 1 0 50324 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_539
timestamp 1666464484
transform 1 0 50692 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1666464484
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_553
timestamp 1666464484
transform 1 0 51980 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_565
timestamp 1666464484
transform 1 0 53084 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_569
timestamp 1666464484
transform 1 0 53452 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_571
timestamp 1666464484
transform 1 0 53636 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_583
timestamp 1666464484
transform 1 0 54740 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_595
timestamp 1666464484
transform 1 0 55844 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_599
timestamp 1666464484
transform 1 0 56212 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_601
timestamp 1666464484
transform 1 0 56396 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_613
timestamp 1666464484
transform 1 0 57500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1666464484
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_16
timestamp 1666464484
transform 1 0 2576 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_28
timestamp 1666464484
transform 1 0 3680 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_40
timestamp 1666464484
transform 1 0 4784 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_44
timestamp 1666464484
transform 1 0 5152 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_46
timestamp 1666464484
transform 1 0 5336 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_58
timestamp 1666464484
transform 1 0 6440 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_70
timestamp 1666464484
transform 1 0 7544 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_74
timestamp 1666464484
transform 1 0 7912 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_76
timestamp 1666464484
transform 1 0 8096 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_88
timestamp 1666464484
transform 1 0 9200 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_100
timestamp 1666464484
transform 1 0 10304 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_104
timestamp 1666464484
transform 1 0 10672 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_106
timestamp 1666464484
transform 1 0 10856 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_118
timestamp 1666464484
transform 1 0 11960 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_130
timestamp 1666464484
transform 1 0 13064 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_134
timestamp 1666464484
transform 1 0 13432 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_136
timestamp 1666464484
transform 1 0 13616 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_148
timestamp 1666464484
transform 1 0 14720 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_160
timestamp 1666464484
transform 1 0 15824 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_164
timestamp 1666464484
transform 1 0 16192 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_166
timestamp 1666464484
transform 1 0 16376 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_178
timestamp 1666464484
transform 1 0 17480 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_190
timestamp 1666464484
transform 1 0 18584 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_194
timestamp 1666464484
transform 1 0 18952 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_196
timestamp 1666464484
transform 1 0 19136 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_208
timestamp 1666464484
transform 1 0 20240 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_220
timestamp 1666464484
transform 1 0 21344 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_224
timestamp 1666464484
transform 1 0 21712 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_226
timestamp 1666464484
transform 1 0 21896 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_238
timestamp 1666464484
transform 1 0 23000 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_250
timestamp 1666464484
transform 1 0 24104 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_254
timestamp 1666464484
transform 1 0 24472 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_256
timestamp 1666464484
transform 1 0 24656 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_268
timestamp 1666464484
transform 1 0 25760 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_280
timestamp 1666464484
transform 1 0 26864 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_284
timestamp 1666464484
transform 1 0 27232 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_286
timestamp 1666464484
transform 1 0 27416 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_298
timestamp 1666464484
transform 1 0 28520 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_310
timestamp 1666464484
transform 1 0 29624 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_314
timestamp 1666464484
transform 1 0 29992 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_316
timestamp 1666464484
transform 1 0 30176 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_328
timestamp 1666464484
transform 1 0 31280 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_340
timestamp 1666464484
transform 1 0 32384 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_344
timestamp 1666464484
transform 1 0 32752 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_346
timestamp 1666464484
transform 1 0 32936 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_358
timestamp 1666464484
transform 1 0 34040 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_370
timestamp 1666464484
transform 1 0 35144 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_374
timestamp 1666464484
transform 1 0 35512 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_376
timestamp 1666464484
transform 1 0 35696 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_388
timestamp 1666464484
transform 1 0 36800 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_400
timestamp 1666464484
transform 1 0 37904 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_404
timestamp 1666464484
transform 1 0 38272 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_406
timestamp 1666464484
transform 1 0 38456 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_418
timestamp 1666464484
transform 1 0 39560 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_430
timestamp 1666464484
transform 1 0 40664 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_434
timestamp 1666464484
transform 1 0 41032 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_436
timestamp 1666464484
transform 1 0 41216 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_448
timestamp 1666464484
transform 1 0 42320 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_460
timestamp 1666464484
transform 1 0 43424 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_464
timestamp 1666464484
transform 1 0 43792 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_466
timestamp 1666464484
transform 1 0 43976 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_478
timestamp 1666464484
transform 1 0 45080 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_490
timestamp 1666464484
transform 1 0 46184 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_494
timestamp 1666464484
transform 1 0 46552 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_496
timestamp 1666464484
transform 1 0 46736 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_508
timestamp 1666464484
transform 1 0 47840 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_520
timestamp 1666464484
transform 1 0 48944 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_524
timestamp 1666464484
transform 1 0 49312 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_526
timestamp 1666464484
transform 1 0 49496 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_538
timestamp 1666464484
transform 1 0 50600 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_550
timestamp 1666464484
transform 1 0 51704 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_554
timestamp 1666464484
transform 1 0 52072 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_556
timestamp 1666464484
transform 1 0 52256 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_568
timestamp 1666464484
transform 1 0 53360 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_580
timestamp 1666464484
transform 1 0 54464 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_584
timestamp 1666464484
transform 1 0 54832 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_586
timestamp 1666464484
transform 1 0 55016 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_598
timestamp 1666464484
transform 1 0 56120 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_610
timestamp 1666464484
transform 1 0 57224 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_614
timestamp 1666464484
transform 1 0 57592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_616
timestamp 1666464484
transform 1 0 57776 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_624
timestamp 1666464484
transform 1 0 58512 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1666464484
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1666464484
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_27
timestamp 1666464484
transform 1 0 3588 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_31
timestamp 1666464484
transform 1 0 3956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_43
timestamp 1666464484
transform 1 0 5060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_55
timestamp 1666464484
transform 1 0 6164 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_59
timestamp 1666464484
transform 1 0 6532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_61
timestamp 1666464484
transform 1 0 6716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_73
timestamp 1666464484
transform 1 0 7820 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_85
timestamp 1666464484
transform 1 0 8924 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_89
timestamp 1666464484
transform 1 0 9292 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_91
timestamp 1666464484
transform 1 0 9476 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_103
timestamp 1666464484
transform 1 0 10580 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_115
timestamp 1666464484
transform 1 0 11684 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_119
timestamp 1666464484
transform 1 0 12052 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_121
timestamp 1666464484
transform 1 0 12236 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_133
timestamp 1666464484
transform 1 0 13340 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_145
timestamp 1666464484
transform 1 0 14444 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_149
timestamp 1666464484
transform 1 0 14812 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_151
timestamp 1666464484
transform 1 0 14996 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_163
timestamp 1666464484
transform 1 0 16100 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_175
timestamp 1666464484
transform 1 0 17204 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_179
timestamp 1666464484
transform 1 0 17572 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1666464484
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1666464484
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_205
timestamp 1666464484
transform 1 0 19964 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_209
timestamp 1666464484
transform 1 0 20332 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_211
timestamp 1666464484
transform 1 0 20516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_223
timestamp 1666464484
transform 1 0 21620 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_235
timestamp 1666464484
transform 1 0 22724 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_239
timestamp 1666464484
transform 1 0 23092 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_241
timestamp 1666464484
transform 1 0 23276 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_253
timestamp 1666464484
transform 1 0 24380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_265
timestamp 1666464484
transform 1 0 25484 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_269
timestamp 1666464484
transform 1 0 25852 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_271
timestamp 1666464484
transform 1 0 26036 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_283
timestamp 1666464484
transform 1 0 27140 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_295
timestamp 1666464484
transform 1 0 28244 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_299
timestamp 1666464484
transform 1 0 28612 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_301
timestamp 1666464484
transform 1 0 28796 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_313
timestamp 1666464484
transform 1 0 29900 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_325
timestamp 1666464484
transform 1 0 31004 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_329
timestamp 1666464484
transform 1 0 31372 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_331
timestamp 1666464484
transform 1 0 31556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_343
timestamp 1666464484
transform 1 0 32660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_355
timestamp 1666464484
transform 1 0 33764 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_359
timestamp 1666464484
transform 1 0 34132 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1666464484
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1666464484
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_385
timestamp 1666464484
transform 1 0 36524 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_389
timestamp 1666464484
transform 1 0 36892 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_391
timestamp 1666464484
transform 1 0 37076 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_403
timestamp 1666464484
transform 1 0 38180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_415
timestamp 1666464484
transform 1 0 39284 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_419
timestamp 1666464484
transform 1 0 39652 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_421
timestamp 1666464484
transform 1 0 39836 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_433
timestamp 1666464484
transform 1 0 40940 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_445
timestamp 1666464484
transform 1 0 42044 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_449
timestamp 1666464484
transform 1 0 42412 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_451
timestamp 1666464484
transform 1 0 42596 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_463
timestamp 1666464484
transform 1 0 43700 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_475
timestamp 1666464484
transform 1 0 44804 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_479
timestamp 1666464484
transform 1 0 45172 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_481
timestamp 1666464484
transform 1 0 45356 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_493
timestamp 1666464484
transform 1 0 46460 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_505
timestamp 1666464484
transform 1 0 47564 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_509
timestamp 1666464484
transform 1 0 47932 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_511
timestamp 1666464484
transform 1 0 48116 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_523
timestamp 1666464484
transform 1 0 49220 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_535
timestamp 1666464484
transform 1 0 50324 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_539
timestamp 1666464484
transform 1 0 50692 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1666464484
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_553
timestamp 1666464484
transform 1 0 51980 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_565
timestamp 1666464484
transform 1 0 53084 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_569
timestamp 1666464484
transform 1 0 53452 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_571
timestamp 1666464484
transform 1 0 53636 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_583
timestamp 1666464484
transform 1 0 54740 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_595
timestamp 1666464484
transform 1 0 55844 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_599
timestamp 1666464484
transform 1 0 56212 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_601
timestamp 1666464484
transform 1 0 56396 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_613
timestamp 1666464484
transform 1 0 57500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1666464484
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_16
timestamp 1666464484
transform 1 0 2576 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_28
timestamp 1666464484
transform 1 0 3680 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_40
timestamp 1666464484
transform 1 0 4784 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_44
timestamp 1666464484
transform 1 0 5152 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_46
timestamp 1666464484
transform 1 0 5336 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_58
timestamp 1666464484
transform 1 0 6440 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_70
timestamp 1666464484
transform 1 0 7544 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_74
timestamp 1666464484
transform 1 0 7912 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_76
timestamp 1666464484
transform 1 0 8096 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_88
timestamp 1666464484
transform 1 0 9200 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_100
timestamp 1666464484
transform 1 0 10304 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_104
timestamp 1666464484
transform 1 0 10672 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_106
timestamp 1666464484
transform 1 0 10856 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_118
timestamp 1666464484
transform 1 0 11960 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_130
timestamp 1666464484
transform 1 0 13064 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_134
timestamp 1666464484
transform 1 0 13432 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_136
timestamp 1666464484
transform 1 0 13616 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_148
timestamp 1666464484
transform 1 0 14720 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_160
timestamp 1666464484
transform 1 0 15824 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_164
timestamp 1666464484
transform 1 0 16192 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_166
timestamp 1666464484
transform 1 0 16376 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_178
timestamp 1666464484
transform 1 0 17480 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_190
timestamp 1666464484
transform 1 0 18584 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_194
timestamp 1666464484
transform 1 0 18952 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_196
timestamp 1666464484
transform 1 0 19136 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_208
timestamp 1666464484
transform 1 0 20240 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_220
timestamp 1666464484
transform 1 0 21344 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_224
timestamp 1666464484
transform 1 0 21712 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_226
timestamp 1666464484
transform 1 0 21896 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_238
timestamp 1666464484
transform 1 0 23000 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_250
timestamp 1666464484
transform 1 0 24104 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_254
timestamp 1666464484
transform 1 0 24472 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_256
timestamp 1666464484
transform 1 0 24656 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_268
timestamp 1666464484
transform 1 0 25760 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_280
timestamp 1666464484
transform 1 0 26864 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_284
timestamp 1666464484
transform 1 0 27232 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_286
timestamp 1666464484
transform 1 0 27416 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_298
timestamp 1666464484
transform 1 0 28520 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_310
timestamp 1666464484
transform 1 0 29624 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_314
timestamp 1666464484
transform 1 0 29992 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_316
timestamp 1666464484
transform 1 0 30176 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_328
timestamp 1666464484
transform 1 0 31280 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_340
timestamp 1666464484
transform 1 0 32384 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_344
timestamp 1666464484
transform 1 0 32752 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_346
timestamp 1666464484
transform 1 0 32936 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_358
timestamp 1666464484
transform 1 0 34040 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_370
timestamp 1666464484
transform 1 0 35144 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_374
timestamp 1666464484
transform 1 0 35512 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_376
timestamp 1666464484
transform 1 0 35696 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_388
timestamp 1666464484
transform 1 0 36800 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_400
timestamp 1666464484
transform 1 0 37904 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_404
timestamp 1666464484
transform 1 0 38272 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_406
timestamp 1666464484
transform 1 0 38456 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_418
timestamp 1666464484
transform 1 0 39560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_430
timestamp 1666464484
transform 1 0 40664 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_434
timestamp 1666464484
transform 1 0 41032 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_436
timestamp 1666464484
transform 1 0 41216 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_448
timestamp 1666464484
transform 1 0 42320 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_460
timestamp 1666464484
transform 1 0 43424 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_464
timestamp 1666464484
transform 1 0 43792 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_466
timestamp 1666464484
transform 1 0 43976 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_478
timestamp 1666464484
transform 1 0 45080 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_490
timestamp 1666464484
transform 1 0 46184 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_494
timestamp 1666464484
transform 1 0 46552 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_496
timestamp 1666464484
transform 1 0 46736 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_508
timestamp 1666464484
transform 1 0 47840 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_520
timestamp 1666464484
transform 1 0 48944 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_524
timestamp 1666464484
transform 1 0 49312 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_526
timestamp 1666464484
transform 1 0 49496 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_538
timestamp 1666464484
transform 1 0 50600 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_550
timestamp 1666464484
transform 1 0 51704 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_554
timestamp 1666464484
transform 1 0 52072 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_556
timestamp 1666464484
transform 1 0 52256 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_568
timestamp 1666464484
transform 1 0 53360 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_580
timestamp 1666464484
transform 1 0 54464 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_584
timestamp 1666464484
transform 1 0 54832 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_586
timestamp 1666464484
transform 1 0 55016 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_598
timestamp 1666464484
transform 1 0 56120 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_610
timestamp 1666464484
transform 1 0 57224 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_614
timestamp 1666464484
transform 1 0 57592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_616
timestamp 1666464484
transform 1 0 57776 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_624
timestamp 1666464484
transform 1 0 58512 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1666464484
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1666464484
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_27
timestamp 1666464484
transform 1 0 3588 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_31
timestamp 1666464484
transform 1 0 3956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_43
timestamp 1666464484
transform 1 0 5060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_55
timestamp 1666464484
transform 1 0 6164 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_59
timestamp 1666464484
transform 1 0 6532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_61
timestamp 1666464484
transform 1 0 6716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_73
timestamp 1666464484
transform 1 0 7820 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_85
timestamp 1666464484
transform 1 0 8924 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_89
timestamp 1666464484
transform 1 0 9292 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_91
timestamp 1666464484
transform 1 0 9476 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_103
timestamp 1666464484
transform 1 0 10580 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_115
timestamp 1666464484
transform 1 0 11684 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_119
timestamp 1666464484
transform 1 0 12052 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_121
timestamp 1666464484
transform 1 0 12236 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_133
timestamp 1666464484
transform 1 0 13340 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_145
timestamp 1666464484
transform 1 0 14444 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_149
timestamp 1666464484
transform 1 0 14812 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_151
timestamp 1666464484
transform 1 0 14996 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_163
timestamp 1666464484
transform 1 0 16100 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_175
timestamp 1666464484
transform 1 0 17204 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_179
timestamp 1666464484
transform 1 0 17572 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1666464484
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1666464484
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_205
timestamp 1666464484
transform 1 0 19964 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_209
timestamp 1666464484
transform 1 0 20332 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_211
timestamp 1666464484
transform 1 0 20516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_223
timestamp 1666464484
transform 1 0 21620 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_235
timestamp 1666464484
transform 1 0 22724 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_239
timestamp 1666464484
transform 1 0 23092 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_241
timestamp 1666464484
transform 1 0 23276 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_253
timestamp 1666464484
transform 1 0 24380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_265
timestamp 1666464484
transform 1 0 25484 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_269
timestamp 1666464484
transform 1 0 25852 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_271
timestamp 1666464484
transform 1 0 26036 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_283
timestamp 1666464484
transform 1 0 27140 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_295
timestamp 1666464484
transform 1 0 28244 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_299
timestamp 1666464484
transform 1 0 28612 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_301
timestamp 1666464484
transform 1 0 28796 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_313
timestamp 1666464484
transform 1 0 29900 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_325
timestamp 1666464484
transform 1 0 31004 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_329
timestamp 1666464484
transform 1 0 31372 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_331
timestamp 1666464484
transform 1 0 31556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_343
timestamp 1666464484
transform 1 0 32660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_355
timestamp 1666464484
transform 1 0 33764 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_359
timestamp 1666464484
transform 1 0 34132 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1666464484
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1666464484
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_385
timestamp 1666464484
transform 1 0 36524 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_389
timestamp 1666464484
transform 1 0 36892 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_391
timestamp 1666464484
transform 1 0 37076 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_403
timestamp 1666464484
transform 1 0 38180 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_415
timestamp 1666464484
transform 1 0 39284 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_419
timestamp 1666464484
transform 1 0 39652 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_421
timestamp 1666464484
transform 1 0 39836 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_433
timestamp 1666464484
transform 1 0 40940 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_445
timestamp 1666464484
transform 1 0 42044 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_449
timestamp 1666464484
transform 1 0 42412 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_451
timestamp 1666464484
transform 1 0 42596 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_463
timestamp 1666464484
transform 1 0 43700 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_475
timestamp 1666464484
transform 1 0 44804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_479
timestamp 1666464484
transform 1 0 45172 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_481
timestamp 1666464484
transform 1 0 45356 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_493
timestamp 1666464484
transform 1 0 46460 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_505
timestamp 1666464484
transform 1 0 47564 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_509
timestamp 1666464484
transform 1 0 47932 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_511
timestamp 1666464484
transform 1 0 48116 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_523
timestamp 1666464484
transform 1 0 49220 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_535
timestamp 1666464484
transform 1 0 50324 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_539
timestamp 1666464484
transform 1 0 50692 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1666464484
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_553
timestamp 1666464484
transform 1 0 51980 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_565
timestamp 1666464484
transform 1 0 53084 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_569
timestamp 1666464484
transform 1 0 53452 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_571
timestamp 1666464484
transform 1 0 53636 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_583
timestamp 1666464484
transform 1 0 54740 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_595
timestamp 1666464484
transform 1 0 55844 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_599
timestamp 1666464484
transform 1 0 56212 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_601
timestamp 1666464484
transform 1 0 56396 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_613
timestamp 1666464484
transform 1 0 57500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1666464484
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_16
timestamp 1666464484
transform 1 0 2576 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_28
timestamp 1666464484
transform 1 0 3680 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_40
timestamp 1666464484
transform 1 0 4784 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_44
timestamp 1666464484
transform 1 0 5152 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_46
timestamp 1666464484
transform 1 0 5336 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_58
timestamp 1666464484
transform 1 0 6440 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_70
timestamp 1666464484
transform 1 0 7544 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_74
timestamp 1666464484
transform 1 0 7912 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_76
timestamp 1666464484
transform 1 0 8096 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_88
timestamp 1666464484
transform 1 0 9200 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_100
timestamp 1666464484
transform 1 0 10304 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_104
timestamp 1666464484
transform 1 0 10672 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_106
timestamp 1666464484
transform 1 0 10856 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_118
timestamp 1666464484
transform 1 0 11960 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_130
timestamp 1666464484
transform 1 0 13064 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_134
timestamp 1666464484
transform 1 0 13432 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_136
timestamp 1666464484
transform 1 0 13616 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_148
timestamp 1666464484
transform 1 0 14720 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_160
timestamp 1666464484
transform 1 0 15824 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_164
timestamp 1666464484
transform 1 0 16192 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_166
timestamp 1666464484
transform 1 0 16376 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_178
timestamp 1666464484
transform 1 0 17480 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_190
timestamp 1666464484
transform 1 0 18584 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_194
timestamp 1666464484
transform 1 0 18952 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_196
timestamp 1666464484
transform 1 0 19136 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_208
timestamp 1666464484
transform 1 0 20240 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_220
timestamp 1666464484
transform 1 0 21344 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_224
timestamp 1666464484
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_226
timestamp 1666464484
transform 1 0 21896 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_238
timestamp 1666464484
transform 1 0 23000 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_250
timestamp 1666464484
transform 1 0 24104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_254
timestamp 1666464484
transform 1 0 24472 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_256
timestamp 1666464484
transform 1 0 24656 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_268
timestamp 1666464484
transform 1 0 25760 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_280
timestamp 1666464484
transform 1 0 26864 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_284
timestamp 1666464484
transform 1 0 27232 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_286
timestamp 1666464484
transform 1 0 27416 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_298
timestamp 1666464484
transform 1 0 28520 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_310
timestamp 1666464484
transform 1 0 29624 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_314
timestamp 1666464484
transform 1 0 29992 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_316
timestamp 1666464484
transform 1 0 30176 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_328
timestamp 1666464484
transform 1 0 31280 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_340
timestamp 1666464484
transform 1 0 32384 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_344
timestamp 1666464484
transform 1 0 32752 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_346
timestamp 1666464484
transform 1 0 32936 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_358
timestamp 1666464484
transform 1 0 34040 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_370
timestamp 1666464484
transform 1 0 35144 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_374
timestamp 1666464484
transform 1 0 35512 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_376
timestamp 1666464484
transform 1 0 35696 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_388
timestamp 1666464484
transform 1 0 36800 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_400
timestamp 1666464484
transform 1 0 37904 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_404
timestamp 1666464484
transform 1 0 38272 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_406
timestamp 1666464484
transform 1 0 38456 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_418
timestamp 1666464484
transform 1 0 39560 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_430
timestamp 1666464484
transform 1 0 40664 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_434
timestamp 1666464484
transform 1 0 41032 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_436
timestamp 1666464484
transform 1 0 41216 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_448
timestamp 1666464484
transform 1 0 42320 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_460
timestamp 1666464484
transform 1 0 43424 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_464
timestamp 1666464484
transform 1 0 43792 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_466
timestamp 1666464484
transform 1 0 43976 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_478
timestamp 1666464484
transform 1 0 45080 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_490
timestamp 1666464484
transform 1 0 46184 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_494
timestamp 1666464484
transform 1 0 46552 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_496
timestamp 1666464484
transform 1 0 46736 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_508
timestamp 1666464484
transform 1 0 47840 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_520
timestamp 1666464484
transform 1 0 48944 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_524
timestamp 1666464484
transform 1 0 49312 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_526
timestamp 1666464484
transform 1 0 49496 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_538
timestamp 1666464484
transform 1 0 50600 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_550
timestamp 1666464484
transform 1 0 51704 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_554
timestamp 1666464484
transform 1 0 52072 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_556
timestamp 1666464484
transform 1 0 52256 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_568
timestamp 1666464484
transform 1 0 53360 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_580
timestamp 1666464484
transform 1 0 54464 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_584
timestamp 1666464484
transform 1 0 54832 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_586
timestamp 1666464484
transform 1 0 55016 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_598
timestamp 1666464484
transform 1 0 56120 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_610
timestamp 1666464484
transform 1 0 57224 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_614
timestamp 1666464484
transform 1 0 57592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_616
timestamp 1666464484
transform 1 0 57776 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_624
timestamp 1666464484
transform 1 0 58512 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1666464484
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1666464484
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_27
timestamp 1666464484
transform 1 0 3588 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_31
timestamp 1666464484
transform 1 0 3956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_43
timestamp 1666464484
transform 1 0 5060 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_55
timestamp 1666464484
transform 1 0 6164 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_59
timestamp 1666464484
transform 1 0 6532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_61
timestamp 1666464484
transform 1 0 6716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_73
timestamp 1666464484
transform 1 0 7820 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_85
timestamp 1666464484
transform 1 0 8924 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_89
timestamp 1666464484
transform 1 0 9292 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_91
timestamp 1666464484
transform 1 0 9476 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_103
timestamp 1666464484
transform 1 0 10580 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_115
timestamp 1666464484
transform 1 0 11684 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_119
timestamp 1666464484
transform 1 0 12052 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_121
timestamp 1666464484
transform 1 0 12236 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_133
timestamp 1666464484
transform 1 0 13340 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_145
timestamp 1666464484
transform 1 0 14444 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_149
timestamp 1666464484
transform 1 0 14812 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_151
timestamp 1666464484
transform 1 0 14996 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_163
timestamp 1666464484
transform 1 0 16100 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_175
timestamp 1666464484
transform 1 0 17204 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_179
timestamp 1666464484
transform 1 0 17572 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1666464484
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1666464484
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_205
timestamp 1666464484
transform 1 0 19964 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_209
timestamp 1666464484
transform 1 0 20332 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_211
timestamp 1666464484
transform 1 0 20516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_223
timestamp 1666464484
transform 1 0 21620 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_235
timestamp 1666464484
transform 1 0 22724 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_239
timestamp 1666464484
transform 1 0 23092 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_241
timestamp 1666464484
transform 1 0 23276 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_253
timestamp 1666464484
transform 1 0 24380 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_265
timestamp 1666464484
transform 1 0 25484 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_269
timestamp 1666464484
transform 1 0 25852 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_271
timestamp 1666464484
transform 1 0 26036 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_283
timestamp 1666464484
transform 1 0 27140 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_295
timestamp 1666464484
transform 1 0 28244 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_299
timestamp 1666464484
transform 1 0 28612 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_301
timestamp 1666464484
transform 1 0 28796 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_313
timestamp 1666464484
transform 1 0 29900 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_325
timestamp 1666464484
transform 1 0 31004 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_329
timestamp 1666464484
transform 1 0 31372 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_331
timestamp 1666464484
transform 1 0 31556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_343
timestamp 1666464484
transform 1 0 32660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_355
timestamp 1666464484
transform 1 0 33764 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_359
timestamp 1666464484
transform 1 0 34132 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1666464484
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1666464484
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_385
timestamp 1666464484
transform 1 0 36524 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_389
timestamp 1666464484
transform 1 0 36892 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_391
timestamp 1666464484
transform 1 0 37076 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_403
timestamp 1666464484
transform 1 0 38180 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_415
timestamp 1666464484
transform 1 0 39284 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_419
timestamp 1666464484
transform 1 0 39652 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_421
timestamp 1666464484
transform 1 0 39836 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_433
timestamp 1666464484
transform 1 0 40940 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_445
timestamp 1666464484
transform 1 0 42044 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_449
timestamp 1666464484
transform 1 0 42412 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_451
timestamp 1666464484
transform 1 0 42596 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_463
timestamp 1666464484
transform 1 0 43700 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_475
timestamp 1666464484
transform 1 0 44804 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_479
timestamp 1666464484
transform 1 0 45172 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_481
timestamp 1666464484
transform 1 0 45356 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_493
timestamp 1666464484
transform 1 0 46460 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_505
timestamp 1666464484
transform 1 0 47564 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_509
timestamp 1666464484
transform 1 0 47932 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_511
timestamp 1666464484
transform 1 0 48116 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_523
timestamp 1666464484
transform 1 0 49220 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_535
timestamp 1666464484
transform 1 0 50324 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_539
timestamp 1666464484
transform 1 0 50692 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1666464484
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_553
timestamp 1666464484
transform 1 0 51980 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_565
timestamp 1666464484
transform 1 0 53084 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_569
timestamp 1666464484
transform 1 0 53452 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_571
timestamp 1666464484
transform 1 0 53636 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_583
timestamp 1666464484
transform 1 0 54740 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_595
timestamp 1666464484
transform 1 0 55844 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_599
timestamp 1666464484
transform 1 0 56212 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_601
timestamp 1666464484
transform 1 0 56396 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_613
timestamp 1666464484
transform 1 0 57500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1666464484
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_16
timestamp 1666464484
transform 1 0 2576 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_28
timestamp 1666464484
transform 1 0 3680 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_40
timestamp 1666464484
transform 1 0 4784 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_44
timestamp 1666464484
transform 1 0 5152 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_46
timestamp 1666464484
transform 1 0 5336 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_58
timestamp 1666464484
transform 1 0 6440 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_70
timestamp 1666464484
transform 1 0 7544 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_74
timestamp 1666464484
transform 1 0 7912 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_76
timestamp 1666464484
transform 1 0 8096 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_88
timestamp 1666464484
transform 1 0 9200 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_100
timestamp 1666464484
transform 1 0 10304 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_104
timestamp 1666464484
transform 1 0 10672 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_106
timestamp 1666464484
transform 1 0 10856 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_118
timestamp 1666464484
transform 1 0 11960 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_130
timestamp 1666464484
transform 1 0 13064 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_134
timestamp 1666464484
transform 1 0 13432 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_136
timestamp 1666464484
transform 1 0 13616 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_148
timestamp 1666464484
transform 1 0 14720 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_160
timestamp 1666464484
transform 1 0 15824 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_164
timestamp 1666464484
transform 1 0 16192 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_166
timestamp 1666464484
transform 1 0 16376 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_178
timestamp 1666464484
transform 1 0 17480 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_190
timestamp 1666464484
transform 1 0 18584 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_194
timestamp 1666464484
transform 1 0 18952 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_196
timestamp 1666464484
transform 1 0 19136 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_208
timestamp 1666464484
transform 1 0 20240 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_220
timestamp 1666464484
transform 1 0 21344 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_224
timestamp 1666464484
transform 1 0 21712 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_226
timestamp 1666464484
transform 1 0 21896 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_238
timestamp 1666464484
transform 1 0 23000 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_250
timestamp 1666464484
transform 1 0 24104 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_254
timestamp 1666464484
transform 1 0 24472 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_256
timestamp 1666464484
transform 1 0 24656 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_268
timestamp 1666464484
transform 1 0 25760 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_280
timestamp 1666464484
transform 1 0 26864 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_284
timestamp 1666464484
transform 1 0 27232 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_286
timestamp 1666464484
transform 1 0 27416 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_298
timestamp 1666464484
transform 1 0 28520 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_310
timestamp 1666464484
transform 1 0 29624 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_314
timestamp 1666464484
transform 1 0 29992 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_316
timestamp 1666464484
transform 1 0 30176 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_328
timestamp 1666464484
transform 1 0 31280 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_340
timestamp 1666464484
transform 1 0 32384 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_344
timestamp 1666464484
transform 1 0 32752 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_346
timestamp 1666464484
transform 1 0 32936 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_358
timestamp 1666464484
transform 1 0 34040 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_370
timestamp 1666464484
transform 1 0 35144 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_374
timestamp 1666464484
transform 1 0 35512 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_376
timestamp 1666464484
transform 1 0 35696 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_388
timestamp 1666464484
transform 1 0 36800 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_400
timestamp 1666464484
transform 1 0 37904 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_404
timestamp 1666464484
transform 1 0 38272 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_406
timestamp 1666464484
transform 1 0 38456 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_418
timestamp 1666464484
transform 1 0 39560 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_430
timestamp 1666464484
transform 1 0 40664 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_434
timestamp 1666464484
transform 1 0 41032 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_436
timestamp 1666464484
transform 1 0 41216 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_448
timestamp 1666464484
transform 1 0 42320 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_460
timestamp 1666464484
transform 1 0 43424 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_464
timestamp 1666464484
transform 1 0 43792 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_466
timestamp 1666464484
transform 1 0 43976 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_478
timestamp 1666464484
transform 1 0 45080 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_490
timestamp 1666464484
transform 1 0 46184 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_494
timestamp 1666464484
transform 1 0 46552 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_496
timestamp 1666464484
transform 1 0 46736 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_508
timestamp 1666464484
transform 1 0 47840 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_520
timestamp 1666464484
transform 1 0 48944 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_524
timestamp 1666464484
transform 1 0 49312 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_526
timestamp 1666464484
transform 1 0 49496 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_538
timestamp 1666464484
transform 1 0 50600 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_550
timestamp 1666464484
transform 1 0 51704 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_554
timestamp 1666464484
transform 1 0 52072 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_556
timestamp 1666464484
transform 1 0 52256 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_568
timestamp 1666464484
transform 1 0 53360 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_580
timestamp 1666464484
transform 1 0 54464 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_584
timestamp 1666464484
transform 1 0 54832 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_586
timestamp 1666464484
transform 1 0 55016 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_598
timestamp 1666464484
transform 1 0 56120 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_610
timestamp 1666464484
transform 1 0 57224 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_614
timestamp 1666464484
transform 1 0 57592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_616
timestamp 1666464484
transform 1 0 57776 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_624
timestamp 1666464484
transform 1 0 58512 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1666464484
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1666464484
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_27
timestamp 1666464484
transform 1 0 3588 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_31
timestamp 1666464484
transform 1 0 3956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_43
timestamp 1666464484
transform 1 0 5060 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_55
timestamp 1666464484
transform 1 0 6164 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_59
timestamp 1666464484
transform 1 0 6532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_61
timestamp 1666464484
transform 1 0 6716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_73
timestamp 1666464484
transform 1 0 7820 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_85
timestamp 1666464484
transform 1 0 8924 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_89
timestamp 1666464484
transform 1 0 9292 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_91
timestamp 1666464484
transform 1 0 9476 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_103
timestamp 1666464484
transform 1 0 10580 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_115
timestamp 1666464484
transform 1 0 11684 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_119
timestamp 1666464484
transform 1 0 12052 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_121
timestamp 1666464484
transform 1 0 12236 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_133
timestamp 1666464484
transform 1 0 13340 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_145
timestamp 1666464484
transform 1 0 14444 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_149
timestamp 1666464484
transform 1 0 14812 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_151
timestamp 1666464484
transform 1 0 14996 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_163
timestamp 1666464484
transform 1 0 16100 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_175
timestamp 1666464484
transform 1 0 17204 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_179
timestamp 1666464484
transform 1 0 17572 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1666464484
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1666464484
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_205
timestamp 1666464484
transform 1 0 19964 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_209
timestamp 1666464484
transform 1 0 20332 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_211
timestamp 1666464484
transform 1 0 20516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_223
timestamp 1666464484
transform 1 0 21620 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_235
timestamp 1666464484
transform 1 0 22724 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_239
timestamp 1666464484
transform 1 0 23092 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_241
timestamp 1666464484
transform 1 0 23276 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_253
timestamp 1666464484
transform 1 0 24380 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_265
timestamp 1666464484
transform 1 0 25484 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_269
timestamp 1666464484
transform 1 0 25852 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_271
timestamp 1666464484
transform 1 0 26036 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_283
timestamp 1666464484
transform 1 0 27140 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_295
timestamp 1666464484
transform 1 0 28244 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_299
timestamp 1666464484
transform 1 0 28612 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_301
timestamp 1666464484
transform 1 0 28796 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_313
timestamp 1666464484
transform 1 0 29900 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_325
timestamp 1666464484
transform 1 0 31004 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_329
timestamp 1666464484
transform 1 0 31372 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_331
timestamp 1666464484
transform 1 0 31556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_343
timestamp 1666464484
transform 1 0 32660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_355
timestamp 1666464484
transform 1 0 33764 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_359
timestamp 1666464484
transform 1 0 34132 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1666464484
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1666464484
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_385
timestamp 1666464484
transform 1 0 36524 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_389
timestamp 1666464484
transform 1 0 36892 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_391
timestamp 1666464484
transform 1 0 37076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_403
timestamp 1666464484
transform 1 0 38180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_415
timestamp 1666464484
transform 1 0 39284 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_419
timestamp 1666464484
transform 1 0 39652 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_421
timestamp 1666464484
transform 1 0 39836 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_433
timestamp 1666464484
transform 1 0 40940 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_445
timestamp 1666464484
transform 1 0 42044 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_449
timestamp 1666464484
transform 1 0 42412 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_451
timestamp 1666464484
transform 1 0 42596 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_463
timestamp 1666464484
transform 1 0 43700 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_475
timestamp 1666464484
transform 1 0 44804 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_479
timestamp 1666464484
transform 1 0 45172 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_481
timestamp 1666464484
transform 1 0 45356 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_493
timestamp 1666464484
transform 1 0 46460 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_505
timestamp 1666464484
transform 1 0 47564 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_509
timestamp 1666464484
transform 1 0 47932 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_511
timestamp 1666464484
transform 1 0 48116 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_523
timestamp 1666464484
transform 1 0 49220 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_535
timestamp 1666464484
transform 1 0 50324 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_539
timestamp 1666464484
transform 1 0 50692 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1666464484
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_553
timestamp 1666464484
transform 1 0 51980 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_565
timestamp 1666464484
transform 1 0 53084 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_569
timestamp 1666464484
transform 1 0 53452 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_571
timestamp 1666464484
transform 1 0 53636 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_583
timestamp 1666464484
transform 1 0 54740 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_595
timestamp 1666464484
transform 1 0 55844 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_599
timestamp 1666464484
transform 1 0 56212 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_601
timestamp 1666464484
transform 1 0 56396 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_613
timestamp 1666464484
transform 1 0 57500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1666464484
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_16
timestamp 1666464484
transform 1 0 2576 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_28
timestamp 1666464484
transform 1 0 3680 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_40
timestamp 1666464484
transform 1 0 4784 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_44
timestamp 1666464484
transform 1 0 5152 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_46
timestamp 1666464484
transform 1 0 5336 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_58
timestamp 1666464484
transform 1 0 6440 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_70
timestamp 1666464484
transform 1 0 7544 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_74
timestamp 1666464484
transform 1 0 7912 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_76
timestamp 1666464484
transform 1 0 8096 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_88
timestamp 1666464484
transform 1 0 9200 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_100
timestamp 1666464484
transform 1 0 10304 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_104
timestamp 1666464484
transform 1 0 10672 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_106
timestamp 1666464484
transform 1 0 10856 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_118
timestamp 1666464484
transform 1 0 11960 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_130
timestamp 1666464484
transform 1 0 13064 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_134
timestamp 1666464484
transform 1 0 13432 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_136
timestamp 1666464484
transform 1 0 13616 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_148
timestamp 1666464484
transform 1 0 14720 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_160
timestamp 1666464484
transform 1 0 15824 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_164
timestamp 1666464484
transform 1 0 16192 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_166
timestamp 1666464484
transform 1 0 16376 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_178
timestamp 1666464484
transform 1 0 17480 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_190
timestamp 1666464484
transform 1 0 18584 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_194
timestamp 1666464484
transform 1 0 18952 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_196
timestamp 1666464484
transform 1 0 19136 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_208
timestamp 1666464484
transform 1 0 20240 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_220
timestamp 1666464484
transform 1 0 21344 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_224
timestamp 1666464484
transform 1 0 21712 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_226
timestamp 1666464484
transform 1 0 21896 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_238
timestamp 1666464484
transform 1 0 23000 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_250
timestamp 1666464484
transform 1 0 24104 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_254
timestamp 1666464484
transform 1 0 24472 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_256
timestamp 1666464484
transform 1 0 24656 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_268
timestamp 1666464484
transform 1 0 25760 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_280
timestamp 1666464484
transform 1 0 26864 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_284
timestamp 1666464484
transform 1 0 27232 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_286
timestamp 1666464484
transform 1 0 27416 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_298
timestamp 1666464484
transform 1 0 28520 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_310
timestamp 1666464484
transform 1 0 29624 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_314
timestamp 1666464484
transform 1 0 29992 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_316
timestamp 1666464484
transform 1 0 30176 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_328
timestamp 1666464484
transform 1 0 31280 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_340
timestamp 1666464484
transform 1 0 32384 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_344
timestamp 1666464484
transform 1 0 32752 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_346
timestamp 1666464484
transform 1 0 32936 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_358
timestamp 1666464484
transform 1 0 34040 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_370
timestamp 1666464484
transform 1 0 35144 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_374
timestamp 1666464484
transform 1 0 35512 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_376
timestamp 1666464484
transform 1 0 35696 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_388
timestamp 1666464484
transform 1 0 36800 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_400
timestamp 1666464484
transform 1 0 37904 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_404
timestamp 1666464484
transform 1 0 38272 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_406
timestamp 1666464484
transform 1 0 38456 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_418
timestamp 1666464484
transform 1 0 39560 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_430
timestamp 1666464484
transform 1 0 40664 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_434
timestamp 1666464484
transform 1 0 41032 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_436
timestamp 1666464484
transform 1 0 41216 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_448
timestamp 1666464484
transform 1 0 42320 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_460
timestamp 1666464484
transform 1 0 43424 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_464
timestamp 1666464484
transform 1 0 43792 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_466
timestamp 1666464484
transform 1 0 43976 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_478
timestamp 1666464484
transform 1 0 45080 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_490
timestamp 1666464484
transform 1 0 46184 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_494
timestamp 1666464484
transform 1 0 46552 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_496
timestamp 1666464484
transform 1 0 46736 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_508
timestamp 1666464484
transform 1 0 47840 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_520
timestamp 1666464484
transform 1 0 48944 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_524
timestamp 1666464484
transform 1 0 49312 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_526
timestamp 1666464484
transform 1 0 49496 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_538
timestamp 1666464484
transform 1 0 50600 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_550
timestamp 1666464484
transform 1 0 51704 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_554
timestamp 1666464484
transform 1 0 52072 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_556
timestamp 1666464484
transform 1 0 52256 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_568
timestamp 1666464484
transform 1 0 53360 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_580
timestamp 1666464484
transform 1 0 54464 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_584
timestamp 1666464484
transform 1 0 54832 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_586
timestamp 1666464484
transform 1 0 55016 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_598
timestamp 1666464484
transform 1 0 56120 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_610
timestamp 1666464484
transform 1 0 57224 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_614
timestamp 1666464484
transform 1 0 57592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_616
timestamp 1666464484
transform 1 0 57776 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_624
timestamp 1666464484
transform 1 0 58512 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1666464484
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1666464484
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_27
timestamp 1666464484
transform 1 0 3588 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_31
timestamp 1666464484
transform 1 0 3956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_43
timestamp 1666464484
transform 1 0 5060 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_55
timestamp 1666464484
transform 1 0 6164 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_59
timestamp 1666464484
transform 1 0 6532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_61
timestamp 1666464484
transform 1 0 6716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_73
timestamp 1666464484
transform 1 0 7820 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_85
timestamp 1666464484
transform 1 0 8924 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_89
timestamp 1666464484
transform 1 0 9292 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_91
timestamp 1666464484
transform 1 0 9476 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_103
timestamp 1666464484
transform 1 0 10580 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_115
timestamp 1666464484
transform 1 0 11684 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_119
timestamp 1666464484
transform 1 0 12052 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_121
timestamp 1666464484
transform 1 0 12236 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_133
timestamp 1666464484
transform 1 0 13340 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_145
timestamp 1666464484
transform 1 0 14444 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_149
timestamp 1666464484
transform 1 0 14812 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_151
timestamp 1666464484
transform 1 0 14996 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_163
timestamp 1666464484
transform 1 0 16100 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_175
timestamp 1666464484
transform 1 0 17204 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_179
timestamp 1666464484
transform 1 0 17572 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1666464484
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1666464484
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_205
timestamp 1666464484
transform 1 0 19964 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_209
timestamp 1666464484
transform 1 0 20332 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_211
timestamp 1666464484
transform 1 0 20516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_223
timestamp 1666464484
transform 1 0 21620 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_235
timestamp 1666464484
transform 1 0 22724 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_239
timestamp 1666464484
transform 1 0 23092 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_241
timestamp 1666464484
transform 1 0 23276 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_253
timestamp 1666464484
transform 1 0 24380 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_265
timestamp 1666464484
transform 1 0 25484 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_269
timestamp 1666464484
transform 1 0 25852 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_271
timestamp 1666464484
transform 1 0 26036 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_283
timestamp 1666464484
transform 1 0 27140 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_295
timestamp 1666464484
transform 1 0 28244 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_299
timestamp 1666464484
transform 1 0 28612 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_301
timestamp 1666464484
transform 1 0 28796 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_313
timestamp 1666464484
transform 1 0 29900 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_325
timestamp 1666464484
transform 1 0 31004 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_329
timestamp 1666464484
transform 1 0 31372 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_331
timestamp 1666464484
transform 1 0 31556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_343
timestamp 1666464484
transform 1 0 32660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_355
timestamp 1666464484
transform 1 0 33764 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_359
timestamp 1666464484
transform 1 0 34132 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1666464484
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1666464484
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_385
timestamp 1666464484
transform 1 0 36524 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_389
timestamp 1666464484
transform 1 0 36892 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_391
timestamp 1666464484
transform 1 0 37076 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_403
timestamp 1666464484
transform 1 0 38180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_415
timestamp 1666464484
transform 1 0 39284 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_419
timestamp 1666464484
transform 1 0 39652 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_421
timestamp 1666464484
transform 1 0 39836 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_433
timestamp 1666464484
transform 1 0 40940 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_445
timestamp 1666464484
transform 1 0 42044 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_449
timestamp 1666464484
transform 1 0 42412 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_451
timestamp 1666464484
transform 1 0 42596 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_463
timestamp 1666464484
transform 1 0 43700 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_475
timestamp 1666464484
transform 1 0 44804 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_479
timestamp 1666464484
transform 1 0 45172 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_481
timestamp 1666464484
transform 1 0 45356 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_493
timestamp 1666464484
transform 1 0 46460 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_505
timestamp 1666464484
transform 1 0 47564 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_509
timestamp 1666464484
transform 1 0 47932 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_511
timestamp 1666464484
transform 1 0 48116 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_523
timestamp 1666464484
transform 1 0 49220 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_535
timestamp 1666464484
transform 1 0 50324 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_539
timestamp 1666464484
transform 1 0 50692 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1666464484
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_553
timestamp 1666464484
transform 1 0 51980 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_565
timestamp 1666464484
transform 1 0 53084 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_569
timestamp 1666464484
transform 1 0 53452 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_571
timestamp 1666464484
transform 1 0 53636 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_583
timestamp 1666464484
transform 1 0 54740 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_595
timestamp 1666464484
transform 1 0 55844 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_599
timestamp 1666464484
transform 1 0 56212 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_601
timestamp 1666464484
transform 1 0 56396 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_613
timestamp 1666464484
transform 1 0 57500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1666464484
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_16
timestamp 1666464484
transform 1 0 2576 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_28
timestamp 1666464484
transform 1 0 3680 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_40
timestamp 1666464484
transform 1 0 4784 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_44
timestamp 1666464484
transform 1 0 5152 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_46
timestamp 1666464484
transform 1 0 5336 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_58
timestamp 1666464484
transform 1 0 6440 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_70
timestamp 1666464484
transform 1 0 7544 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_74
timestamp 1666464484
transform 1 0 7912 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_76
timestamp 1666464484
transform 1 0 8096 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_88
timestamp 1666464484
transform 1 0 9200 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_100
timestamp 1666464484
transform 1 0 10304 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_104
timestamp 1666464484
transform 1 0 10672 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_106
timestamp 1666464484
transform 1 0 10856 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_118
timestamp 1666464484
transform 1 0 11960 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_130
timestamp 1666464484
transform 1 0 13064 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_134
timestamp 1666464484
transform 1 0 13432 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_136
timestamp 1666464484
transform 1 0 13616 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_148
timestamp 1666464484
transform 1 0 14720 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_160
timestamp 1666464484
transform 1 0 15824 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_164
timestamp 1666464484
transform 1 0 16192 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_166
timestamp 1666464484
transform 1 0 16376 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_178
timestamp 1666464484
transform 1 0 17480 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_190
timestamp 1666464484
transform 1 0 18584 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_194
timestamp 1666464484
transform 1 0 18952 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_196
timestamp 1666464484
transform 1 0 19136 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_208
timestamp 1666464484
transform 1 0 20240 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_220
timestamp 1666464484
transform 1 0 21344 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_224
timestamp 1666464484
transform 1 0 21712 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_226
timestamp 1666464484
transform 1 0 21896 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_238
timestamp 1666464484
transform 1 0 23000 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_250
timestamp 1666464484
transform 1 0 24104 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_254
timestamp 1666464484
transform 1 0 24472 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_256
timestamp 1666464484
transform 1 0 24656 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_268
timestamp 1666464484
transform 1 0 25760 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_280
timestamp 1666464484
transform 1 0 26864 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_284
timestamp 1666464484
transform 1 0 27232 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_286
timestamp 1666464484
transform 1 0 27416 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_298
timestamp 1666464484
transform 1 0 28520 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_310
timestamp 1666464484
transform 1 0 29624 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_314
timestamp 1666464484
transform 1 0 29992 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_316
timestamp 1666464484
transform 1 0 30176 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_328
timestamp 1666464484
transform 1 0 31280 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_340
timestamp 1666464484
transform 1 0 32384 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_344
timestamp 1666464484
transform 1 0 32752 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_346
timestamp 1666464484
transform 1 0 32936 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_358
timestamp 1666464484
transform 1 0 34040 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_370
timestamp 1666464484
transform 1 0 35144 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_374
timestamp 1666464484
transform 1 0 35512 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_376
timestamp 1666464484
transform 1 0 35696 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_388
timestamp 1666464484
transform 1 0 36800 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_400
timestamp 1666464484
transform 1 0 37904 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_404
timestamp 1666464484
transform 1 0 38272 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_406
timestamp 1666464484
transform 1 0 38456 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_418
timestamp 1666464484
transform 1 0 39560 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_430
timestamp 1666464484
transform 1 0 40664 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_434
timestamp 1666464484
transform 1 0 41032 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_436
timestamp 1666464484
transform 1 0 41216 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_448
timestamp 1666464484
transform 1 0 42320 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_460
timestamp 1666464484
transform 1 0 43424 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_464
timestamp 1666464484
transform 1 0 43792 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_466
timestamp 1666464484
transform 1 0 43976 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_478
timestamp 1666464484
transform 1 0 45080 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_490
timestamp 1666464484
transform 1 0 46184 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_494
timestamp 1666464484
transform 1 0 46552 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_496
timestamp 1666464484
transform 1 0 46736 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_508
timestamp 1666464484
transform 1 0 47840 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_520
timestamp 1666464484
transform 1 0 48944 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_524
timestamp 1666464484
transform 1 0 49312 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_526
timestamp 1666464484
transform 1 0 49496 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_538
timestamp 1666464484
transform 1 0 50600 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_550
timestamp 1666464484
transform 1 0 51704 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_554
timestamp 1666464484
transform 1 0 52072 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_556
timestamp 1666464484
transform 1 0 52256 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_568
timestamp 1666464484
transform 1 0 53360 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_580
timestamp 1666464484
transform 1 0 54464 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_584
timestamp 1666464484
transform 1 0 54832 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_586
timestamp 1666464484
transform 1 0 55016 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_598
timestamp 1666464484
transform 1 0 56120 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_610
timestamp 1666464484
transform 1 0 57224 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_614
timestamp 1666464484
transform 1 0 57592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_616
timestamp 1666464484
transform 1 0 57776 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_624
timestamp 1666464484
transform 1 0 58512 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1666464484
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1666464484
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_27
timestamp 1666464484
transform 1 0 3588 0 -1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_31
timestamp 1666464484
transform 1 0 3956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_43
timestamp 1666464484
transform 1 0 5060 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_55
timestamp 1666464484
transform 1 0 6164 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_59
timestamp 1666464484
transform 1 0 6532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_61
timestamp 1666464484
transform 1 0 6716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_73
timestamp 1666464484
transform 1 0 7820 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_85
timestamp 1666464484
transform 1 0 8924 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_89
timestamp 1666464484
transform 1 0 9292 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_91
timestamp 1666464484
transform 1 0 9476 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_103
timestamp 1666464484
transform 1 0 10580 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_115
timestamp 1666464484
transform 1 0 11684 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_119
timestamp 1666464484
transform 1 0 12052 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_121
timestamp 1666464484
transform 1 0 12236 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_133
timestamp 1666464484
transform 1 0 13340 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_145
timestamp 1666464484
transform 1 0 14444 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_149
timestamp 1666464484
transform 1 0 14812 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_151
timestamp 1666464484
transform 1 0 14996 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_163
timestamp 1666464484
transform 1 0 16100 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_175
timestamp 1666464484
transform 1 0 17204 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_179
timestamp 1666464484
transform 1 0 17572 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1666464484
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1666464484
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_205
timestamp 1666464484
transform 1 0 19964 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_209
timestamp 1666464484
transform 1 0 20332 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_211
timestamp 1666464484
transform 1 0 20516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_223
timestamp 1666464484
transform 1 0 21620 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_235
timestamp 1666464484
transform 1 0 22724 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_239
timestamp 1666464484
transform 1 0 23092 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_241
timestamp 1666464484
transform 1 0 23276 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_253
timestamp 1666464484
transform 1 0 24380 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_265
timestamp 1666464484
transform 1 0 25484 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_269
timestamp 1666464484
transform 1 0 25852 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_271
timestamp 1666464484
transform 1 0 26036 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_283
timestamp 1666464484
transform 1 0 27140 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_295
timestamp 1666464484
transform 1 0 28244 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_299
timestamp 1666464484
transform 1 0 28612 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_301
timestamp 1666464484
transform 1 0 28796 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_313
timestamp 1666464484
transform 1 0 29900 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_325
timestamp 1666464484
transform 1 0 31004 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_329
timestamp 1666464484
transform 1 0 31372 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_331
timestamp 1666464484
transform 1 0 31556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_343
timestamp 1666464484
transform 1 0 32660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_355
timestamp 1666464484
transform 1 0 33764 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_359
timestamp 1666464484
transform 1 0 34132 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1666464484
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1666464484
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_385
timestamp 1666464484
transform 1 0 36524 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_389
timestamp 1666464484
transform 1 0 36892 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_391
timestamp 1666464484
transform 1 0 37076 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_403
timestamp 1666464484
transform 1 0 38180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_415
timestamp 1666464484
transform 1 0 39284 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_419
timestamp 1666464484
transform 1 0 39652 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_421
timestamp 1666464484
transform 1 0 39836 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_433
timestamp 1666464484
transform 1 0 40940 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_445
timestamp 1666464484
transform 1 0 42044 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_449
timestamp 1666464484
transform 1 0 42412 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_451
timestamp 1666464484
transform 1 0 42596 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_463
timestamp 1666464484
transform 1 0 43700 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_475
timestamp 1666464484
transform 1 0 44804 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_479
timestamp 1666464484
transform 1 0 45172 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_481
timestamp 1666464484
transform 1 0 45356 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_493
timestamp 1666464484
transform 1 0 46460 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_505
timestamp 1666464484
transform 1 0 47564 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_509
timestamp 1666464484
transform 1 0 47932 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_511
timestamp 1666464484
transform 1 0 48116 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_523
timestamp 1666464484
transform 1 0 49220 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_535
timestamp 1666464484
transform 1 0 50324 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_539
timestamp 1666464484
transform 1 0 50692 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1666464484
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_553
timestamp 1666464484
transform 1 0 51980 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_565
timestamp 1666464484
transform 1 0 53084 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_569
timestamp 1666464484
transform 1 0 53452 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_571
timestamp 1666464484
transform 1 0 53636 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_583
timestamp 1666464484
transform 1 0 54740 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_595
timestamp 1666464484
transform 1 0 55844 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_599
timestamp 1666464484
transform 1 0 56212 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_601
timestamp 1666464484
transform 1 0 56396 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_613
timestamp 1666464484
transform 1 0 57500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1666464484
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_16
timestamp 1666464484
transform 1 0 2576 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_28
timestamp 1666464484
transform 1 0 3680 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_40
timestamp 1666464484
transform 1 0 4784 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_44
timestamp 1666464484
transform 1 0 5152 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_46
timestamp 1666464484
transform 1 0 5336 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_58
timestamp 1666464484
transform 1 0 6440 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_70
timestamp 1666464484
transform 1 0 7544 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_74
timestamp 1666464484
transform 1 0 7912 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_76
timestamp 1666464484
transform 1 0 8096 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_88
timestamp 1666464484
transform 1 0 9200 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_100
timestamp 1666464484
transform 1 0 10304 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_104
timestamp 1666464484
transform 1 0 10672 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_106
timestamp 1666464484
transform 1 0 10856 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_118
timestamp 1666464484
transform 1 0 11960 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_130
timestamp 1666464484
transform 1 0 13064 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_134
timestamp 1666464484
transform 1 0 13432 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_136
timestamp 1666464484
transform 1 0 13616 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_148
timestamp 1666464484
transform 1 0 14720 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_160
timestamp 1666464484
transform 1 0 15824 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_164
timestamp 1666464484
transform 1 0 16192 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_166
timestamp 1666464484
transform 1 0 16376 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_178
timestamp 1666464484
transform 1 0 17480 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_190
timestamp 1666464484
transform 1 0 18584 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_194
timestamp 1666464484
transform 1 0 18952 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_196
timestamp 1666464484
transform 1 0 19136 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_208
timestamp 1666464484
transform 1 0 20240 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_220
timestamp 1666464484
transform 1 0 21344 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_224
timestamp 1666464484
transform 1 0 21712 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_226
timestamp 1666464484
transform 1 0 21896 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_238
timestamp 1666464484
transform 1 0 23000 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_250
timestamp 1666464484
transform 1 0 24104 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_254
timestamp 1666464484
transform 1 0 24472 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_256
timestamp 1666464484
transform 1 0 24656 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_268
timestamp 1666464484
transform 1 0 25760 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_280
timestamp 1666464484
transform 1 0 26864 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_284
timestamp 1666464484
transform 1 0 27232 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_286
timestamp 1666464484
transform 1 0 27416 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_298
timestamp 1666464484
transform 1 0 28520 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_310
timestamp 1666464484
transform 1 0 29624 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_314
timestamp 1666464484
transform 1 0 29992 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_316
timestamp 1666464484
transform 1 0 30176 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_328
timestamp 1666464484
transform 1 0 31280 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_340
timestamp 1666464484
transform 1 0 32384 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_344
timestamp 1666464484
transform 1 0 32752 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_346
timestamp 1666464484
transform 1 0 32936 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_358
timestamp 1666464484
transform 1 0 34040 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_370
timestamp 1666464484
transform 1 0 35144 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_374
timestamp 1666464484
transform 1 0 35512 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_376
timestamp 1666464484
transform 1 0 35696 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_388
timestamp 1666464484
transform 1 0 36800 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_400
timestamp 1666464484
transform 1 0 37904 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_404
timestamp 1666464484
transform 1 0 38272 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_406
timestamp 1666464484
transform 1 0 38456 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_418
timestamp 1666464484
transform 1 0 39560 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_430
timestamp 1666464484
transform 1 0 40664 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_434
timestamp 1666464484
transform 1 0 41032 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_436
timestamp 1666464484
transform 1 0 41216 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_448
timestamp 1666464484
transform 1 0 42320 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_460
timestamp 1666464484
transform 1 0 43424 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_464
timestamp 1666464484
transform 1 0 43792 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_466
timestamp 1666464484
transform 1 0 43976 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_478
timestamp 1666464484
transform 1 0 45080 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_490
timestamp 1666464484
transform 1 0 46184 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_494
timestamp 1666464484
transform 1 0 46552 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_496
timestamp 1666464484
transform 1 0 46736 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_508
timestamp 1666464484
transform 1 0 47840 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_520
timestamp 1666464484
transform 1 0 48944 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_524
timestamp 1666464484
transform 1 0 49312 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_526
timestamp 1666464484
transform 1 0 49496 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_538
timestamp 1666464484
transform 1 0 50600 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_550
timestamp 1666464484
transform 1 0 51704 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_554
timestamp 1666464484
transform 1 0 52072 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_556
timestamp 1666464484
transform 1 0 52256 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_568
timestamp 1666464484
transform 1 0 53360 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_580
timestamp 1666464484
transform 1 0 54464 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_584
timestamp 1666464484
transform 1 0 54832 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_586
timestamp 1666464484
transform 1 0 55016 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_598
timestamp 1666464484
transform 1 0 56120 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_610
timestamp 1666464484
transform 1 0 57224 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_614
timestamp 1666464484
transform 1 0 57592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_616
timestamp 1666464484
transform 1 0 57776 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_624
timestamp 1666464484
transform 1 0 58512 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1666464484
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1666464484
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_27
timestamp 1666464484
transform 1 0 3588 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_31
timestamp 1666464484
transform 1 0 3956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_43
timestamp 1666464484
transform 1 0 5060 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_55
timestamp 1666464484
transform 1 0 6164 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_59
timestamp 1666464484
transform 1 0 6532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_61
timestamp 1666464484
transform 1 0 6716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_73
timestamp 1666464484
transform 1 0 7820 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_85
timestamp 1666464484
transform 1 0 8924 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_89
timestamp 1666464484
transform 1 0 9292 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_91
timestamp 1666464484
transform 1 0 9476 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_103
timestamp 1666464484
transform 1 0 10580 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_115
timestamp 1666464484
transform 1 0 11684 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_119
timestamp 1666464484
transform 1 0 12052 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_121
timestamp 1666464484
transform 1 0 12236 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_133
timestamp 1666464484
transform 1 0 13340 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_145
timestamp 1666464484
transform 1 0 14444 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_149
timestamp 1666464484
transform 1 0 14812 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_151
timestamp 1666464484
transform 1 0 14996 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_163
timestamp 1666464484
transform 1 0 16100 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_175
timestamp 1666464484
transform 1 0 17204 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_179
timestamp 1666464484
transform 1 0 17572 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1666464484
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1666464484
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_205
timestamp 1666464484
transform 1 0 19964 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_209
timestamp 1666464484
transform 1 0 20332 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_211
timestamp 1666464484
transform 1 0 20516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_223
timestamp 1666464484
transform 1 0 21620 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_235
timestamp 1666464484
transform 1 0 22724 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_239
timestamp 1666464484
transform 1 0 23092 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_241
timestamp 1666464484
transform 1 0 23276 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_253
timestamp 1666464484
transform 1 0 24380 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_265
timestamp 1666464484
transform 1 0 25484 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_269
timestamp 1666464484
transform 1 0 25852 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_271
timestamp 1666464484
transform 1 0 26036 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_283
timestamp 1666464484
transform 1 0 27140 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_295
timestamp 1666464484
transform 1 0 28244 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_299
timestamp 1666464484
transform 1 0 28612 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_301
timestamp 1666464484
transform 1 0 28796 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_313
timestamp 1666464484
transform 1 0 29900 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_325
timestamp 1666464484
transform 1 0 31004 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_329
timestamp 1666464484
transform 1 0 31372 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_331
timestamp 1666464484
transform 1 0 31556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_343
timestamp 1666464484
transform 1 0 32660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_355
timestamp 1666464484
transform 1 0 33764 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_359
timestamp 1666464484
transform 1 0 34132 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1666464484
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1666464484
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_385
timestamp 1666464484
transform 1 0 36524 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_389
timestamp 1666464484
transform 1 0 36892 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_391
timestamp 1666464484
transform 1 0 37076 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_403
timestamp 1666464484
transform 1 0 38180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_415
timestamp 1666464484
transform 1 0 39284 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_419
timestamp 1666464484
transform 1 0 39652 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_421
timestamp 1666464484
transform 1 0 39836 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_433
timestamp 1666464484
transform 1 0 40940 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_445
timestamp 1666464484
transform 1 0 42044 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_449
timestamp 1666464484
transform 1 0 42412 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_451
timestamp 1666464484
transform 1 0 42596 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_463
timestamp 1666464484
transform 1 0 43700 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_475
timestamp 1666464484
transform 1 0 44804 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_479
timestamp 1666464484
transform 1 0 45172 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_481
timestamp 1666464484
transform 1 0 45356 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_493
timestamp 1666464484
transform 1 0 46460 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_505
timestamp 1666464484
transform 1 0 47564 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_509
timestamp 1666464484
transform 1 0 47932 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_511
timestamp 1666464484
transform 1 0 48116 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_523
timestamp 1666464484
transform 1 0 49220 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_535
timestamp 1666464484
transform 1 0 50324 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_539
timestamp 1666464484
transform 1 0 50692 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1666464484
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_553
timestamp 1666464484
transform 1 0 51980 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_565
timestamp 1666464484
transform 1 0 53084 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_569
timestamp 1666464484
transform 1 0 53452 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_571
timestamp 1666464484
transform 1 0 53636 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_583
timestamp 1666464484
transform 1 0 54740 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_595
timestamp 1666464484
transform 1 0 55844 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_599
timestamp 1666464484
transform 1 0 56212 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_601
timestamp 1666464484
transform 1 0 56396 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_613
timestamp 1666464484
transform 1 0 57500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1666464484
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_16
timestamp 1666464484
transform 1 0 2576 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_28
timestamp 1666464484
transform 1 0 3680 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_40
timestamp 1666464484
transform 1 0 4784 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_44
timestamp 1666464484
transform 1 0 5152 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_46
timestamp 1666464484
transform 1 0 5336 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_58
timestamp 1666464484
transform 1 0 6440 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_70
timestamp 1666464484
transform 1 0 7544 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_74
timestamp 1666464484
transform 1 0 7912 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_76
timestamp 1666464484
transform 1 0 8096 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_88
timestamp 1666464484
transform 1 0 9200 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_100
timestamp 1666464484
transform 1 0 10304 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_104
timestamp 1666464484
transform 1 0 10672 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_106
timestamp 1666464484
transform 1 0 10856 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_118
timestamp 1666464484
transform 1 0 11960 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_130
timestamp 1666464484
transform 1 0 13064 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_134
timestamp 1666464484
transform 1 0 13432 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_136
timestamp 1666464484
transform 1 0 13616 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_148
timestamp 1666464484
transform 1 0 14720 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_160
timestamp 1666464484
transform 1 0 15824 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_164
timestamp 1666464484
transform 1 0 16192 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_166
timestamp 1666464484
transform 1 0 16376 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_178
timestamp 1666464484
transform 1 0 17480 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_190
timestamp 1666464484
transform 1 0 18584 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_194
timestamp 1666464484
transform 1 0 18952 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_196
timestamp 1666464484
transform 1 0 19136 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_208
timestamp 1666464484
transform 1 0 20240 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_220
timestamp 1666464484
transform 1 0 21344 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_224
timestamp 1666464484
transform 1 0 21712 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_226
timestamp 1666464484
transform 1 0 21896 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_238
timestamp 1666464484
transform 1 0 23000 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_250
timestamp 1666464484
transform 1 0 24104 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_254
timestamp 1666464484
transform 1 0 24472 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_256
timestamp 1666464484
transform 1 0 24656 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_268
timestamp 1666464484
transform 1 0 25760 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_280
timestamp 1666464484
transform 1 0 26864 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_284
timestamp 1666464484
transform 1 0 27232 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_286
timestamp 1666464484
transform 1 0 27416 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_298
timestamp 1666464484
transform 1 0 28520 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_310
timestamp 1666464484
transform 1 0 29624 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_314
timestamp 1666464484
transform 1 0 29992 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_316
timestamp 1666464484
transform 1 0 30176 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_328
timestamp 1666464484
transform 1 0 31280 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_340
timestamp 1666464484
transform 1 0 32384 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_344
timestamp 1666464484
transform 1 0 32752 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_346
timestamp 1666464484
transform 1 0 32936 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_358
timestamp 1666464484
transform 1 0 34040 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_366
timestamp 1666464484
transform 1 0 34776 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_371
timestamp 1666464484
transform 1 0 35236 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_376
timestamp 1666464484
transform 1 0 35696 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_388
timestamp 1666464484
transform 1 0 36800 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_400
timestamp 1666464484
transform 1 0 37904 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_404
timestamp 1666464484
transform 1 0 38272 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_406
timestamp 1666464484
transform 1 0 38456 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_418
timestamp 1666464484
transform 1 0 39560 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_430
timestamp 1666464484
transform 1 0 40664 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_434
timestamp 1666464484
transform 1 0 41032 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_436
timestamp 1666464484
transform 1 0 41216 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_448
timestamp 1666464484
transform 1 0 42320 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_460
timestamp 1666464484
transform 1 0 43424 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_464
timestamp 1666464484
transform 1 0 43792 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_466
timestamp 1666464484
transform 1 0 43976 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_478
timestamp 1666464484
transform 1 0 45080 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_490
timestamp 1666464484
transform 1 0 46184 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_494
timestamp 1666464484
transform 1 0 46552 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_496
timestamp 1666464484
transform 1 0 46736 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_508
timestamp 1666464484
transform 1 0 47840 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_520
timestamp 1666464484
transform 1 0 48944 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_524
timestamp 1666464484
transform 1 0 49312 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_526
timestamp 1666464484
transform 1 0 49496 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_538
timestamp 1666464484
transform 1 0 50600 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_550
timestamp 1666464484
transform 1 0 51704 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_554
timestamp 1666464484
transform 1 0 52072 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_556
timestamp 1666464484
transform 1 0 52256 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_568
timestamp 1666464484
transform 1 0 53360 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_580
timestamp 1666464484
transform 1 0 54464 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_584
timestamp 1666464484
transform 1 0 54832 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_586
timestamp 1666464484
transform 1 0 55016 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_598
timestamp 1666464484
transform 1 0 56120 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_610
timestamp 1666464484
transform 1 0 57224 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_614
timestamp 1666464484
transform 1 0 57592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_616
timestamp 1666464484
transform 1 0 57776 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_624
timestamp 1666464484
transform 1 0 58512 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1666464484
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1666464484
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_27
timestamp 1666464484
transform 1 0 3588 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_31
timestamp 1666464484
transform 1 0 3956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_43
timestamp 1666464484
transform 1 0 5060 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_55
timestamp 1666464484
transform 1 0 6164 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_59
timestamp 1666464484
transform 1 0 6532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_61
timestamp 1666464484
transform 1 0 6716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_73
timestamp 1666464484
transform 1 0 7820 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_85
timestamp 1666464484
transform 1 0 8924 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_89
timestamp 1666464484
transform 1 0 9292 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_91
timestamp 1666464484
transform 1 0 9476 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_103
timestamp 1666464484
transform 1 0 10580 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_115
timestamp 1666464484
transform 1 0 11684 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_119
timestamp 1666464484
transform 1 0 12052 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_121
timestamp 1666464484
transform 1 0 12236 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_133
timestamp 1666464484
transform 1 0 13340 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_145
timestamp 1666464484
transform 1 0 14444 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_149
timestamp 1666464484
transform 1 0 14812 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_151
timestamp 1666464484
transform 1 0 14996 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_163
timestamp 1666464484
transform 1 0 16100 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_175
timestamp 1666464484
transform 1 0 17204 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_179
timestamp 1666464484
transform 1 0 17572 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1666464484
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1666464484
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_205
timestamp 1666464484
transform 1 0 19964 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_209
timestamp 1666464484
transform 1 0 20332 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_211
timestamp 1666464484
transform 1 0 20516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_223
timestamp 1666464484
transform 1 0 21620 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_235
timestamp 1666464484
transform 1 0 22724 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_239
timestamp 1666464484
transform 1 0 23092 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_241
timestamp 1666464484
transform 1 0 23276 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_253
timestamp 1666464484
transform 1 0 24380 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_265
timestamp 1666464484
transform 1 0 25484 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_269
timestamp 1666464484
transform 1 0 25852 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_271
timestamp 1666464484
transform 1 0 26036 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_283
timestamp 1666464484
transform 1 0 27140 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_295
timestamp 1666464484
transform 1 0 28244 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_299
timestamp 1666464484
transform 1 0 28612 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_301
timestamp 1666464484
transform 1 0 28796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_305
timestamp 1666464484
transform 1 0 29164 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_308
timestamp 1666464484
transform 1 0 29440 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_312
timestamp 1666464484
transform 1 0 29808 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_315
timestamp 1666464484
transform 1 0 30084 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_93_321
timestamp 1666464484
transform 1 0 30636 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_329
timestamp 1666464484
transform 1 0 31372 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_331
timestamp 1666464484
transform 1 0 31556 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_339
timestamp 1666464484
transform 1 0 32292 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_343
timestamp 1666464484
transform 1 0 32660 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_351
timestamp 1666464484
transform 1 0 33396 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_358
timestamp 1666464484
transform 1 0 34040 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_361
timestamp 1666464484
transform 1 0 34316 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_384
timestamp 1666464484
transform 1 0 36432 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_391
timestamp 1666464484
transform 1 0 37076 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_403
timestamp 1666464484
transform 1 0 38180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_415
timestamp 1666464484
transform 1 0 39284 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_419
timestamp 1666464484
transform 1 0 39652 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_421
timestamp 1666464484
transform 1 0 39836 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_429
timestamp 1666464484
transform 1 0 40572 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_432
timestamp 1666464484
transform 1 0 40848 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_444
timestamp 1666464484
transform 1 0 41952 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_451
timestamp 1666464484
transform 1 0 42596 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_463
timestamp 1666464484
transform 1 0 43700 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_475
timestamp 1666464484
transform 1 0 44804 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_479
timestamp 1666464484
transform 1 0 45172 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_481
timestamp 1666464484
transform 1 0 45356 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_493
timestamp 1666464484
transform 1 0 46460 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_505
timestamp 1666464484
transform 1 0 47564 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_509
timestamp 1666464484
transform 1 0 47932 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_511
timestamp 1666464484
transform 1 0 48116 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_523
timestamp 1666464484
transform 1 0 49220 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_535
timestamp 1666464484
transform 1 0 50324 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_539
timestamp 1666464484
transform 1 0 50692 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1666464484
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_553
timestamp 1666464484
transform 1 0 51980 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_565
timestamp 1666464484
transform 1 0 53084 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_569
timestamp 1666464484
transform 1 0 53452 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_571
timestamp 1666464484
transform 1 0 53636 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_583
timestamp 1666464484
transform 1 0 54740 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_595
timestamp 1666464484
transform 1 0 55844 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_599
timestamp 1666464484
transform 1 0 56212 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_601
timestamp 1666464484
transform 1 0 56396 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_613
timestamp 1666464484
transform 1 0 57500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1666464484
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_16
timestamp 1666464484
transform 1 0 2576 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_28
timestamp 1666464484
transform 1 0 3680 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_40
timestamp 1666464484
transform 1 0 4784 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_44
timestamp 1666464484
transform 1 0 5152 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_46
timestamp 1666464484
transform 1 0 5336 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_58
timestamp 1666464484
transform 1 0 6440 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_70
timestamp 1666464484
transform 1 0 7544 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_74
timestamp 1666464484
transform 1 0 7912 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_76
timestamp 1666464484
transform 1 0 8096 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_88
timestamp 1666464484
transform 1 0 9200 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_100
timestamp 1666464484
transform 1 0 10304 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_104
timestamp 1666464484
transform 1 0 10672 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_106
timestamp 1666464484
transform 1 0 10856 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_118
timestamp 1666464484
transform 1 0 11960 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_130
timestamp 1666464484
transform 1 0 13064 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_134
timestamp 1666464484
transform 1 0 13432 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_136
timestamp 1666464484
transform 1 0 13616 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_148
timestamp 1666464484
transform 1 0 14720 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_160
timestamp 1666464484
transform 1 0 15824 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_164
timestamp 1666464484
transform 1 0 16192 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_166
timestamp 1666464484
transform 1 0 16376 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_178
timestamp 1666464484
transform 1 0 17480 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_190
timestamp 1666464484
transform 1 0 18584 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_194
timestamp 1666464484
transform 1 0 18952 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_196
timestamp 1666464484
transform 1 0 19136 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_208
timestamp 1666464484
transform 1 0 20240 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_220
timestamp 1666464484
transform 1 0 21344 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_224
timestamp 1666464484
transform 1 0 21712 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_226
timestamp 1666464484
transform 1 0 21896 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_238
timestamp 1666464484
transform 1 0 23000 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_250
timestamp 1666464484
transform 1 0 24104 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_254
timestamp 1666464484
transform 1 0 24472 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_256
timestamp 1666464484
transform 1 0 24656 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_268
timestamp 1666464484
transform 1 0 25760 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_280
timestamp 1666464484
transform 1 0 26864 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_284
timestamp 1666464484
transform 1 0 27232 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_286
timestamp 1666464484
transform 1 0 27416 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_94_294
timestamp 1666464484
transform 1 0 28152 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_300
timestamp 1666464484
transform 1 0 28704 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_306
timestamp 1666464484
transform 1 0 29256 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_311
timestamp 1666464484
transform 1 0 29716 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_316
timestamp 1666464484
transform 1 0 30176 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_321
timestamp 1666464484
transform 1 0 30636 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_325
timestamp 1666464484
transform 1 0 31004 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_328
timestamp 1666464484
transform 1 0 31280 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_334
timestamp 1666464484
transform 1 0 31832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_337
timestamp 1666464484
transform 1 0 32108 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_343
timestamp 1666464484
transform 1 0 32660 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_346
timestamp 1666464484
transform 1 0 32936 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_353
timestamp 1666464484
transform 1 0 33580 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_359
timestamp 1666464484
transform 1 0 34132 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_365
timestamp 1666464484
transform 1 0 34684 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_371
timestamp 1666464484
transform 1 0 35236 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_376
timestamp 1666464484
transform 1 0 35696 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_380
timestamp 1666464484
transform 1 0 36064 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_386
timestamp 1666464484
transform 1 0 36616 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_392
timestamp 1666464484
transform 1 0 37168 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_398
timestamp 1666464484
transform 1 0 37720 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_404
timestamp 1666464484
transform 1 0 38272 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_406
timestamp 1666464484
transform 1 0 38456 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_410
timestamp 1666464484
transform 1 0 38824 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_414
timestamp 1666464484
transform 1 0 39192 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_417
timestamp 1666464484
transform 1 0 39468 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_423
timestamp 1666464484
transform 1 0 40020 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_429
timestamp 1666464484
transform 1 0 40572 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_94_436
timestamp 1666464484
transform 1 0 41216 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_440
timestamp 1666464484
transform 1 0 41584 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_446
timestamp 1666464484
transform 1 0 42136 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_458
timestamp 1666464484
transform 1 0 43240 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_464
timestamp 1666464484
transform 1 0 43792 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_466
timestamp 1666464484
transform 1 0 43976 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_478
timestamp 1666464484
transform 1 0 45080 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_490
timestamp 1666464484
transform 1 0 46184 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_494
timestamp 1666464484
transform 1 0 46552 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_496
timestamp 1666464484
transform 1 0 46736 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_508
timestamp 1666464484
transform 1 0 47840 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_520
timestamp 1666464484
transform 1 0 48944 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_524
timestamp 1666464484
transform 1 0 49312 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_526
timestamp 1666464484
transform 1 0 49496 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_538
timestamp 1666464484
transform 1 0 50600 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_550
timestamp 1666464484
transform 1 0 51704 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_554
timestamp 1666464484
transform 1 0 52072 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_556
timestamp 1666464484
transform 1 0 52256 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_568
timestamp 1666464484
transform 1 0 53360 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_580
timestamp 1666464484
transform 1 0 54464 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_584
timestamp 1666464484
transform 1 0 54832 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_586
timestamp 1666464484
transform 1 0 55016 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_598
timestamp 1666464484
transform 1 0 56120 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_610
timestamp 1666464484
transform 1 0 57224 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_614
timestamp 1666464484
transform 1 0 57592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_616
timestamp 1666464484
transform 1 0 57776 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_624
timestamp 1666464484
transform 1 0 58512 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1666464484
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1666464484
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_27
timestamp 1666464484
transform 1 0 3588 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_31
timestamp 1666464484
transform 1 0 3956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_43
timestamp 1666464484
transform 1 0 5060 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_55
timestamp 1666464484
transform 1 0 6164 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_59
timestamp 1666464484
transform 1 0 6532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_61
timestamp 1666464484
transform 1 0 6716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_73
timestamp 1666464484
transform 1 0 7820 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_85
timestamp 1666464484
transform 1 0 8924 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_89
timestamp 1666464484
transform 1 0 9292 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_91
timestamp 1666464484
transform 1 0 9476 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_103
timestamp 1666464484
transform 1 0 10580 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_115
timestamp 1666464484
transform 1 0 11684 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_119
timestamp 1666464484
transform 1 0 12052 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_121
timestamp 1666464484
transform 1 0 12236 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_133
timestamp 1666464484
transform 1 0 13340 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_145
timestamp 1666464484
transform 1 0 14444 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_149
timestamp 1666464484
transform 1 0 14812 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_151
timestamp 1666464484
transform 1 0 14996 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_163
timestamp 1666464484
transform 1 0 16100 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_175
timestamp 1666464484
transform 1 0 17204 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_179
timestamp 1666464484
transform 1 0 17572 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1666464484
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1666464484
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_205
timestamp 1666464484
transform 1 0 19964 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_209
timestamp 1666464484
transform 1 0 20332 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_211
timestamp 1666464484
transform 1 0 20516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_223
timestamp 1666464484
transform 1 0 21620 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_235
timestamp 1666464484
transform 1 0 22724 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_239
timestamp 1666464484
transform 1 0 23092 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_241
timestamp 1666464484
transform 1 0 23276 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_253
timestamp 1666464484
transform 1 0 24380 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_265
timestamp 1666464484
transform 1 0 25484 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_269
timestamp 1666464484
transform 1 0 25852 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_271
timestamp 1666464484
transform 1 0 26036 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_275
timestamp 1666464484
transform 1 0 26404 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_282
timestamp 1666464484
transform 1 0 27048 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_288
timestamp 1666464484
transform 1 0 27600 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_291
timestamp 1666464484
transform 1 0 27876 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_298
timestamp 1666464484
transform 1 0 28520 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_301
timestamp 1666464484
transform 1 0 28796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_310
timestamp 1666464484
transform 1 0 29624 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_319
timestamp 1666464484
transform 1 0 30452 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_326
timestamp 1666464484
transform 1 0 31096 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_331
timestamp 1666464484
transform 1 0 31556 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_341
timestamp 1666464484
transform 1 0 32476 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_351
timestamp 1666464484
transform 1 0 33396 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_358
timestamp 1666464484
transform 1 0 34040 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_361
timestamp 1666464484
transform 1 0 34316 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_369
timestamp 1666464484
transform 1 0 35052 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_376
timestamp 1666464484
transform 1 0 35696 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_382
timestamp 1666464484
transform 1 0 36248 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_388
timestamp 1666464484
transform 1 0 36800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_391
timestamp 1666464484
transform 1 0 37076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_396
timestamp 1666464484
transform 1 0 37536 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_403
timestamp 1666464484
transform 1 0 38180 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_410
timestamp 1666464484
transform 1 0 38824 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_414
timestamp 1666464484
transform 1 0 39192 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_418
timestamp 1666464484
transform 1 0 39560 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_421
timestamp 1666464484
transform 1 0 39836 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_427
timestamp 1666464484
transform 1 0 40388 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_431
timestamp 1666464484
transform 1 0 40756 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_438
timestamp 1666464484
transform 1 0 41400 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_95_447
timestamp 1666464484
transform 1 0 42228 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_451
timestamp 1666464484
transform 1 0 42596 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_455
timestamp 1666464484
transform 1 0 42964 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_95_465
timestamp 1666464484
transform 1 0 43884 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_477
timestamp 1666464484
transform 1 0 44988 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_481
timestamp 1666464484
transform 1 0 45356 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_493
timestamp 1666464484
transform 1 0 46460 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_505
timestamp 1666464484
transform 1 0 47564 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_509
timestamp 1666464484
transform 1 0 47932 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_511
timestamp 1666464484
transform 1 0 48116 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_523
timestamp 1666464484
transform 1 0 49220 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_535
timestamp 1666464484
transform 1 0 50324 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_539
timestamp 1666464484
transform 1 0 50692 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1666464484
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_553
timestamp 1666464484
transform 1 0 51980 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_565
timestamp 1666464484
transform 1 0 53084 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_569
timestamp 1666464484
transform 1 0 53452 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_571
timestamp 1666464484
transform 1 0 53636 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_583
timestamp 1666464484
transform 1 0 54740 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_595
timestamp 1666464484
transform 1 0 55844 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_599
timestamp 1666464484
transform 1 0 56212 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_601
timestamp 1666464484
transform 1 0 56396 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_613
timestamp 1666464484
transform 1 0 57500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1666464484
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_16
timestamp 1666464484
transform 1 0 2576 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_28
timestamp 1666464484
transform 1 0 3680 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_40
timestamp 1666464484
transform 1 0 4784 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_44
timestamp 1666464484
transform 1 0 5152 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_46
timestamp 1666464484
transform 1 0 5336 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_58
timestamp 1666464484
transform 1 0 6440 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_70
timestamp 1666464484
transform 1 0 7544 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_74
timestamp 1666464484
transform 1 0 7912 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_76
timestamp 1666464484
transform 1 0 8096 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_88
timestamp 1666464484
transform 1 0 9200 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_100
timestamp 1666464484
transform 1 0 10304 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_104
timestamp 1666464484
transform 1 0 10672 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_106
timestamp 1666464484
transform 1 0 10856 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_118
timestamp 1666464484
transform 1 0 11960 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_130
timestamp 1666464484
transform 1 0 13064 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_134
timestamp 1666464484
transform 1 0 13432 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_136
timestamp 1666464484
transform 1 0 13616 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_148
timestamp 1666464484
transform 1 0 14720 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_160
timestamp 1666464484
transform 1 0 15824 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_164
timestamp 1666464484
transform 1 0 16192 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_166
timestamp 1666464484
transform 1 0 16376 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_178
timestamp 1666464484
transform 1 0 17480 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_190
timestamp 1666464484
transform 1 0 18584 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_194
timestamp 1666464484
transform 1 0 18952 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_196
timestamp 1666464484
transform 1 0 19136 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_208
timestamp 1666464484
transform 1 0 20240 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_220
timestamp 1666464484
transform 1 0 21344 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_224
timestamp 1666464484
transform 1 0 21712 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_226
timestamp 1666464484
transform 1 0 21896 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_238
timestamp 1666464484
transform 1 0 23000 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_250
timestamp 1666464484
transform 1 0 24104 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_254
timestamp 1666464484
transform 1 0 24472 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_256
timestamp 1666464484
transform 1 0 24656 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_262
timestamp 1666464484
transform 1 0 25208 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_269
timestamp 1666464484
transform 1 0 25852 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_273
timestamp 1666464484
transform 1 0 26220 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_276
timestamp 1666464484
transform 1 0 26496 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_283
timestamp 1666464484
transform 1 0 27140 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_96_286
timestamp 1666464484
transform 1 0 27416 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_96_295
timestamp 1666464484
transform 1 0 28244 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_306
timestamp 1666464484
transform 1 0 29256 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_313
timestamp 1666464484
transform 1 0 29900 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_316
timestamp 1666464484
transform 1 0 30176 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_325
timestamp 1666464484
transform 1 0 31004 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_332
timestamp 1666464484
transform 1 0 31648 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_343
timestamp 1666464484
transform 1 0 32660 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_96_346
timestamp 1666464484
transform 1 0 32936 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_352
timestamp 1666464484
transform 1 0 33488 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_361
timestamp 1666464484
transform 1 0 34316 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_96_372
timestamp 1666464484
transform 1 0 35328 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_376
timestamp 1666464484
transform 1 0 35696 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_384
timestamp 1666464484
transform 1 0 36432 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_391
timestamp 1666464484
transform 1 0 37076 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_397
timestamp 1666464484
transform 1 0 37628 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_403
timestamp 1666464484
transform 1 0 38180 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_406
timestamp 1666464484
transform 1 0 38456 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_413
timestamp 1666464484
transform 1 0 39100 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_422
timestamp 1666464484
transform 1 0 39928 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_96_432
timestamp 1666464484
transform 1 0 40848 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_436
timestamp 1666464484
transform 1 0 41216 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_96_445
timestamp 1666464484
transform 1 0 42044 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_451
timestamp 1666464484
transform 1 0 42596 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_456
timestamp 1666464484
transform 1 0 43056 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_463
timestamp 1666464484
transform 1 0 43700 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_96_466
timestamp 1666464484
transform 1 0 43976 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_474
timestamp 1666464484
transform 1 0 44712 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_486
timestamp 1666464484
transform 1 0 45816 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_494
timestamp 1666464484
transform 1 0 46552 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_496
timestamp 1666464484
transform 1 0 46736 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_508
timestamp 1666464484
transform 1 0 47840 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_520
timestamp 1666464484
transform 1 0 48944 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_524
timestamp 1666464484
transform 1 0 49312 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_526
timestamp 1666464484
transform 1 0 49496 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_538
timestamp 1666464484
transform 1 0 50600 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_550
timestamp 1666464484
transform 1 0 51704 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_554
timestamp 1666464484
transform 1 0 52072 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_556
timestamp 1666464484
transform 1 0 52256 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_568
timestamp 1666464484
transform 1 0 53360 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_580
timestamp 1666464484
transform 1 0 54464 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_584
timestamp 1666464484
transform 1 0 54832 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_586
timestamp 1666464484
transform 1 0 55016 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_598
timestamp 1666464484
transform 1 0 56120 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_610
timestamp 1666464484
transform 1 0 57224 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_614
timestamp 1666464484
transform 1 0 57592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_616
timestamp 1666464484
transform 1 0 57776 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_624
timestamp 1666464484
transform 1 0 58512 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1666464484
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1666464484
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_27
timestamp 1666464484
transform 1 0 3588 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_31
timestamp 1666464484
transform 1 0 3956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_43
timestamp 1666464484
transform 1 0 5060 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_55
timestamp 1666464484
transform 1 0 6164 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_59
timestamp 1666464484
transform 1 0 6532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_61
timestamp 1666464484
transform 1 0 6716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_73
timestamp 1666464484
transform 1 0 7820 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_85
timestamp 1666464484
transform 1 0 8924 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_89
timestamp 1666464484
transform 1 0 9292 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_91
timestamp 1666464484
transform 1 0 9476 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_103
timestamp 1666464484
transform 1 0 10580 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_115
timestamp 1666464484
transform 1 0 11684 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_119
timestamp 1666464484
transform 1 0 12052 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_121
timestamp 1666464484
transform 1 0 12236 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_133
timestamp 1666464484
transform 1 0 13340 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_145
timestamp 1666464484
transform 1 0 14444 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_149
timestamp 1666464484
transform 1 0 14812 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_151
timestamp 1666464484
transform 1 0 14996 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_163
timestamp 1666464484
transform 1 0 16100 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_175
timestamp 1666464484
transform 1 0 17204 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_179
timestamp 1666464484
transform 1 0 17572 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1666464484
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1666464484
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_205
timestamp 1666464484
transform 1 0 19964 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_209
timestamp 1666464484
transform 1 0 20332 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_211
timestamp 1666464484
transform 1 0 20516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_223
timestamp 1666464484
transform 1 0 21620 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_235
timestamp 1666464484
transform 1 0 22724 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_239
timestamp 1666464484
transform 1 0 23092 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_241
timestamp 1666464484
transform 1 0 23276 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_97_252
timestamp 1666464484
transform 1 0 24288 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_97_261
timestamp 1666464484
transform 1 0 25116 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_268
timestamp 1666464484
transform 1 0 25760 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_271
timestamp 1666464484
transform 1 0 26036 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_278
timestamp 1666464484
transform 1 0 26680 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_97_286
timestamp 1666464484
transform 1 0 27416 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_97_298
timestamp 1666464484
transform 1 0 28520 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_97_301
timestamp 1666464484
transform 1 0 28796 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_311
timestamp 1666464484
transform 1 0 29716 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_319
timestamp 1666464484
transform 1 0 30452 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_328
timestamp 1666464484
transform 1 0 31280 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_97_331
timestamp 1666464484
transform 1 0 31556 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_340
timestamp 1666464484
transform 1 0 32384 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_350
timestamp 1666464484
transform 1 0 33304 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_97_357
timestamp 1666464484
transform 1 0 33948 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_361
timestamp 1666464484
transform 1 0 34316 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_370
timestamp 1666464484
transform 1 0 35144 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_377
timestamp 1666464484
transform 1 0 35788 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_97_384
timestamp 1666464484
transform 1 0 36432 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_97_391
timestamp 1666464484
transform 1 0 37076 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_396
timestamp 1666464484
transform 1 0 37536 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_400
timestamp 1666464484
transform 1 0 37904 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_406
timestamp 1666464484
transform 1 0 38456 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_97_417
timestamp 1666464484
transform 1 0 39468 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_421
timestamp 1666464484
transform 1 0 39836 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_431
timestamp 1666464484
transform 1 0 40756 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_439
timestamp 1666464484
transform 1 0 41492 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_448
timestamp 1666464484
transform 1 0 42320 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_451
timestamp 1666464484
transform 1 0 42596 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_460
timestamp 1666464484
transform 1 0 43424 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_470
timestamp 1666464484
transform 1 0 44344 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_97_477
timestamp 1666464484
transform 1 0 44988 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_481
timestamp 1666464484
transform 1 0 45356 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_485
timestamp 1666464484
transform 1 0 45724 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_491
timestamp 1666464484
transform 1 0 46276 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_503
timestamp 1666464484
transform 1 0 47380 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_509
timestamp 1666464484
transform 1 0 47932 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_511
timestamp 1666464484
transform 1 0 48116 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_523
timestamp 1666464484
transform 1 0 49220 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_535
timestamp 1666464484
transform 1 0 50324 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_539
timestamp 1666464484
transform 1 0 50692 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1666464484
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_553
timestamp 1666464484
transform 1 0 51980 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_565
timestamp 1666464484
transform 1 0 53084 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_569
timestamp 1666464484
transform 1 0 53452 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_571
timestamp 1666464484
transform 1 0 53636 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_583
timestamp 1666464484
transform 1 0 54740 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_595
timestamp 1666464484
transform 1 0 55844 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_599
timestamp 1666464484
transform 1 0 56212 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_601
timestamp 1666464484
transform 1 0 56396 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_613
timestamp 1666464484
transform 1 0 57500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1666464484
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_16
timestamp 1666464484
transform 1 0 2576 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_28
timestamp 1666464484
transform 1 0 3680 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_40
timestamp 1666464484
transform 1 0 4784 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_44
timestamp 1666464484
transform 1 0 5152 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_46
timestamp 1666464484
transform 1 0 5336 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_58
timestamp 1666464484
transform 1 0 6440 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_70
timestamp 1666464484
transform 1 0 7544 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_74
timestamp 1666464484
transform 1 0 7912 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_76
timestamp 1666464484
transform 1 0 8096 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_88
timestamp 1666464484
transform 1 0 9200 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_100
timestamp 1666464484
transform 1 0 10304 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_104
timestamp 1666464484
transform 1 0 10672 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_106
timestamp 1666464484
transform 1 0 10856 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_118
timestamp 1666464484
transform 1 0 11960 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_130
timestamp 1666464484
transform 1 0 13064 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_134
timestamp 1666464484
transform 1 0 13432 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_136
timestamp 1666464484
transform 1 0 13616 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_148
timestamp 1666464484
transform 1 0 14720 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_160
timestamp 1666464484
transform 1 0 15824 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_164
timestamp 1666464484
transform 1 0 16192 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_166
timestamp 1666464484
transform 1 0 16376 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_178
timestamp 1666464484
transform 1 0 17480 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_190
timestamp 1666464484
transform 1 0 18584 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_194
timestamp 1666464484
transform 1 0 18952 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_196
timestamp 1666464484
transform 1 0 19136 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_208
timestamp 1666464484
transform 1 0 20240 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_220
timestamp 1666464484
transform 1 0 21344 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_224
timestamp 1666464484
transform 1 0 21712 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_226
timestamp 1666464484
transform 1 0 21896 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_240
timestamp 1666464484
transform 1 0 23184 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_246
timestamp 1666464484
transform 1 0 23736 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_253
timestamp 1666464484
transform 1 0 24380 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_98_256
timestamp 1666464484
transform 1 0 24656 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_98_265
timestamp 1666464484
transform 1 0 25484 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_273
timestamp 1666464484
transform 1 0 26220 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_98_283
timestamp 1666464484
transform 1 0 27140 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_286
timestamp 1666464484
transform 1 0 27416 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_295
timestamp 1666464484
transform 1 0 28244 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_306
timestamp 1666464484
transform 1 0 29256 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_313
timestamp 1666464484
transform 1 0 29900 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_98_316
timestamp 1666464484
transform 1 0 30176 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_322
timestamp 1666464484
transform 1 0 30728 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_331
timestamp 1666464484
transform 1 0 31556 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_341
timestamp 1666464484
transform 1 0 32476 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_346
timestamp 1666464484
transform 1 0 32936 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_98_353
timestamp 1666464484
transform 1 0 33580 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_98_366
timestamp 1666464484
transform 1 0 34776 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_373
timestamp 1666464484
transform 1 0 35420 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_376
timestamp 1666464484
transform 1 0 35696 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_383
timestamp 1666464484
transform 1 0 36340 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_387
timestamp 1666464484
transform 1 0 36708 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_393
timestamp 1666464484
transform 1 0 37260 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_403
timestamp 1666464484
transform 1 0 38180 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_406
timestamp 1666464484
transform 1 0 38456 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_98_415
timestamp 1666464484
transform 1 0 39284 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_98_429
timestamp 1666464484
transform 1 0 40572 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_98_436
timestamp 1666464484
transform 1 0 41216 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_444
timestamp 1666464484
transform 1 0 41952 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_454
timestamp 1666464484
transform 1 0 42872 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_463
timestamp 1666464484
transform 1 0 43700 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_466
timestamp 1666464484
transform 1 0 43976 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_473
timestamp 1666464484
transform 1 0 44620 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_480
timestamp 1666464484
transform 1 0 45264 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_487
timestamp 1666464484
transform 1 0 45908 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_493
timestamp 1666464484
transform 1 0 46460 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_496
timestamp 1666464484
transform 1 0 46736 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_98_500
timestamp 1666464484
transform 1 0 47104 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_98_510
timestamp 1666464484
transform 1 0 48024 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_522
timestamp 1666464484
transform 1 0 49128 0 1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_98_526
timestamp 1666464484
transform 1 0 49496 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_538
timestamp 1666464484
transform 1 0 50600 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_550
timestamp 1666464484
transform 1 0 51704 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_554
timestamp 1666464484
transform 1 0 52072 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_556
timestamp 1666464484
transform 1 0 52256 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_568
timestamp 1666464484
transform 1 0 53360 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_580
timestamp 1666464484
transform 1 0 54464 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_584
timestamp 1666464484
transform 1 0 54832 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_586
timestamp 1666464484
transform 1 0 55016 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_598
timestamp 1666464484
transform 1 0 56120 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_610
timestamp 1666464484
transform 1 0 57224 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_614
timestamp 1666464484
transform 1 0 57592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_616
timestamp 1666464484
transform 1 0 57776 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_624
timestamp 1666464484
transform 1 0 58512 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1666464484
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1666464484
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_27
timestamp 1666464484
transform 1 0 3588 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_99_31
timestamp 1666464484
transform 1 0 3956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_43
timestamp 1666464484
transform 1 0 5060 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_55
timestamp 1666464484
transform 1 0 6164 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_59
timestamp 1666464484
transform 1 0 6532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_61
timestamp 1666464484
transform 1 0 6716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_73
timestamp 1666464484
transform 1 0 7820 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_85
timestamp 1666464484
transform 1 0 8924 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_89
timestamp 1666464484
transform 1 0 9292 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_91
timestamp 1666464484
transform 1 0 9476 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_103
timestamp 1666464484
transform 1 0 10580 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_115
timestamp 1666464484
transform 1 0 11684 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_119
timestamp 1666464484
transform 1 0 12052 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_121
timestamp 1666464484
transform 1 0 12236 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_133
timestamp 1666464484
transform 1 0 13340 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_145
timestamp 1666464484
transform 1 0 14444 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_149
timestamp 1666464484
transform 1 0 14812 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_151
timestamp 1666464484
transform 1 0 14996 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_163
timestamp 1666464484
transform 1 0 16100 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_175
timestamp 1666464484
transform 1 0 17204 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_179
timestamp 1666464484
transform 1 0 17572 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1666464484
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1666464484
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_205
timestamp 1666464484
transform 1 0 19964 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_209
timestamp 1666464484
transform 1 0 20332 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_211
timestamp 1666464484
transform 1 0 20516 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_223
timestamp 1666464484
transform 1 0 21620 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_231
timestamp 1666464484
transform 1 0 22356 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_99_237
timestamp 1666464484
transform 1 0 22908 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_241
timestamp 1666464484
transform 1 0 23276 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_245
timestamp 1666464484
transform 1 0 23644 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_254
timestamp 1666464484
transform 1 0 24472 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_262
timestamp 1666464484
transform 1 0 25208 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_268
timestamp 1666464484
transform 1 0 25760 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_271
timestamp 1666464484
transform 1 0 26036 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_279
timestamp 1666464484
transform 1 0 26772 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_288
timestamp 1666464484
transform 1 0 27600 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_292
timestamp 1666464484
transform 1 0 27968 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_298
timestamp 1666464484
transform 1 0 28520 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_301
timestamp 1666464484
transform 1 0 28796 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_311
timestamp 1666464484
transform 1 0 29716 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_320
timestamp 1666464484
transform 1 0 30544 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_99_327
timestamp 1666464484
transform 1 0 31188 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_331
timestamp 1666464484
transform 1 0 31556 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_339
timestamp 1666464484
transform 1 0 32292 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_349
timestamp 1666464484
transform 1 0 33212 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_353
timestamp 1666464484
transform 1 0 33580 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_358
timestamp 1666464484
transform 1 0 34040 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_361
timestamp 1666464484
transform 1 0 34316 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_367
timestamp 1666464484
transform 1 0 34868 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_379
timestamp 1666464484
transform 1 0 35972 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_388
timestamp 1666464484
transform 1 0 36800 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_391
timestamp 1666464484
transform 1 0 37076 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_400
timestamp 1666464484
transform 1 0 37904 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_410
timestamp 1666464484
transform 1 0 38824 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_418
timestamp 1666464484
transform 1 0 39560 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_421
timestamp 1666464484
transform 1 0 39836 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_431
timestamp 1666464484
transform 1 0 40756 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_441
timestamp 1666464484
transform 1 0 41676 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_448
timestamp 1666464484
transform 1 0 42320 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_451
timestamp 1666464484
transform 1 0 42596 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_460
timestamp 1666464484
transform 1 0 43424 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_471
timestamp 1666464484
transform 1 0 44436 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_478
timestamp 1666464484
transform 1 0 45080 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_481
timestamp 1666464484
transform 1 0 45356 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_486
timestamp 1666464484
transform 1 0 45816 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_493
timestamp 1666464484
transform 1 0 46460 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_500
timestamp 1666464484
transform 1 0 47104 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_99_507
timestamp 1666464484
transform 1 0 47748 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_511
timestamp 1666464484
transform 1 0 48116 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_99_516
timestamp 1666464484
transform 1 0 48576 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_522
timestamp 1666464484
transform 1 0 49128 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_525
timestamp 1666464484
transform 1 0 49404 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_537
timestamp 1666464484
transform 1 0 50508 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_541
timestamp 1666464484
transform 1 0 50876 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_545
timestamp 1666464484
transform 1 0 51244 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_551
timestamp 1666464484
transform 1 0 51796 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_99_559
timestamp 1666464484
transform 1 0 52532 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_567
timestamp 1666464484
transform 1 0 53268 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_571
timestamp 1666464484
transform 1 0 53636 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_575
timestamp 1666464484
transform 1 0 54004 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_589
timestamp 1666464484
transform 1 0 55292 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_597
timestamp 1666464484
transform 1 0 56028 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_99_601
timestamp 1666464484
transform 1 0 56396 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_613
timestamp 1666464484
transform 1 0 57500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1666464484
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_16
timestamp 1666464484
transform 1 0 2576 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_28
timestamp 1666464484
transform 1 0 3680 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_36
timestamp 1666464484
transform 1 0 4416 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_100_42
timestamp 1666464484
transform 1 0 4968 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_100_46
timestamp 1666464484
transform 1 0 5336 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_100_55
timestamp 1666464484
transform 1 0 6164 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_62
timestamp 1666464484
transform 1 0 6808 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_74
timestamp 1666464484
transform 1 0 7912 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_76
timestamp 1666464484
transform 1 0 8096 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_87
timestamp 1666464484
transform 1 0 9108 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_102
timestamp 1666464484
transform 1 0 10488 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_100_106
timestamp 1666464484
transform 1 0 10856 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_117
timestamp 1666464484
transform 1 0 11868 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_132
timestamp 1666464484
transform 1 0 13248 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_100_136
timestamp 1666464484
transform 1 0 13616 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_147
timestamp 1666464484
transform 1 0 14628 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_162
timestamp 1666464484
transform 1 0 16008 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_100_166
timestamp 1666464484
transform 1 0 16376 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1666464484
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_192
timestamp 1666464484
transform 1 0 18768 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_100_196
timestamp 1666464484
transform 1 0 19136 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_207
timestamp 1666464484
transform 1 0 20148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_222
timestamp 1666464484
transform 1 0 21528 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_226
timestamp 1666464484
transform 1 0 21896 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_233
timestamp 1666464484
transform 1 0 22540 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_241
timestamp 1666464484
transform 1 0 23276 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_253
timestamp 1666464484
transform 1 0 24380 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_256
timestamp 1666464484
transform 1 0 24656 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_260
timestamp 1666464484
transform 1 0 25024 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_269
timestamp 1666464484
transform 1 0 25852 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_100_283
timestamp 1666464484
transform 1 0 27140 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_286
timestamp 1666464484
transform 1 0 27416 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_100_295
timestamp 1666464484
transform 1 0 28244 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_303
timestamp 1666464484
transform 1 0 28980 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_313
timestamp 1666464484
transform 1 0 29900 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_100_316
timestamp 1666464484
transform 1 0 30176 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_100_329
timestamp 1666464484
transform 1 0 31372 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_341
timestamp 1666464484
transform 1 0 32476 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_100_346
timestamp 1666464484
transform 1 0 32936 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_356
timestamp 1666464484
transform 1 0 33856 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_366
timestamp 1666464484
transform 1 0 34776 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_373
timestamp 1666464484
transform 1 0 35420 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_100_376
timestamp 1666464484
transform 1 0 35696 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_389
timestamp 1666464484
transform 1 0 36892 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_399
timestamp 1666464484
transform 1 0 37812 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_100_406
timestamp 1666464484
transform 1 0 38456 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_415
timestamp 1666464484
transform 1 0 39284 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_421
timestamp 1666464484
transform 1 0 39836 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_433
timestamp 1666464484
transform 1 0 40940 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_100_436
timestamp 1666464484
transform 1 0 41216 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_446
timestamp 1666464484
transform 1 0 42136 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_456
timestamp 1666464484
transform 1 0 43056 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_463
timestamp 1666464484
transform 1 0 43700 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_466
timestamp 1666464484
transform 1 0 43976 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_478
timestamp 1666464484
transform 1 0 45080 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_485
timestamp 1666464484
transform 1 0 45724 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_100_492
timestamp 1666464484
transform 1 0 46368 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_100_496
timestamp 1666464484
transform 1 0 46736 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_501
timestamp 1666464484
transform 1 0 47196 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_508
timestamp 1666464484
transform 1 0 47840 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_515
timestamp 1666464484
transform 1 0 48484 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_100_522
timestamp 1666464484
transform 1 0 49128 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_100_526
timestamp 1666464484
transform 1 0 49496 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_531
timestamp 1666464484
transform 1 0 49956 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_538
timestamp 1666464484
transform 1 0 50600 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_545
timestamp 1666464484
transform 1 0 51244 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_100_552
timestamp 1666464484
transform 1 0 51888 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_100_556
timestamp 1666464484
transform 1 0 52256 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_561
timestamp 1666464484
transform 1 0 52716 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_568
timestamp 1666464484
transform 1 0 53360 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_575
timestamp 1666464484
transform 1 0 54004 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_100_582
timestamp 1666464484
transform 1 0 54648 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_100_586
timestamp 1666464484
transform 1 0 55016 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_100_591
timestamp 1666464484
transform 1 0 55476 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_602
timestamp 1666464484
transform 1 0 56488 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_614
timestamp 1666464484
transform 1 0 57592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_616
timestamp 1666464484
transform 1 0 57776 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_624
timestamp 1666464484
transform 1 0 58512 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1666464484
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_16
timestamp 1666464484
transform 1 0 2576 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_24
timestamp 1666464484
transform 1 0 3312 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_28
timestamp 1666464484
transform 1 0 3680 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_31
timestamp 1666464484
transform 1 0 3956 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_37
timestamp 1666464484
transform 1 0 4508 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_46
timestamp 1666464484
transform 1 0 5336 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_52
timestamp 1666464484
transform 1 0 5888 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_58
timestamp 1666464484
transform 1 0 6440 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_61
timestamp 1666464484
transform 1 0 6716 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_72
timestamp 1666464484
transform 1 0 7728 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_76
timestamp 1666464484
transform 1 0 8096 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_81
timestamp 1666464484
transform 1 0 8556 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_88
timestamp 1666464484
transform 1 0 9200 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_91
timestamp 1666464484
transform 1 0 9476 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_103
timestamp 1666464484
transform 1 0 10580 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_106
timestamp 1666464484
transform 1 0 10856 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_110
timestamp 1666464484
transform 1 0 11224 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_118
timestamp 1666464484
transform 1 0 11960 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_121
timestamp 1666464484
transform 1 0 12236 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_133
timestamp 1666464484
transform 1 0 13340 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_136
timestamp 1666464484
transform 1 0 13616 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_148
timestamp 1666464484
transform 1 0 14720 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_151
timestamp 1666464484
transform 1 0 14996 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_163
timestamp 1666464484
transform 1 0 16100 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_166
timestamp 1666464484
transform 1 0 16376 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_178
timestamp 1666464484
transform 1 0 17480 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_181
timestamp 1666464484
transform 1 0 17756 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_193
timestamp 1666464484
transform 1 0 18860 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_196
timestamp 1666464484
transform 1 0 19136 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_208
timestamp 1666464484
transform 1 0 20240 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_211
timestamp 1666464484
transform 1 0 20516 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_215
timestamp 1666464484
transform 1 0 20884 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_223
timestamp 1666464484
transform 1 0 21620 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_226
timestamp 1666464484
transform 1 0 21896 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_230
timestamp 1666464484
transform 1 0 22264 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_238
timestamp 1666464484
transform 1 0 23000 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_241
timestamp 1666464484
transform 1 0 23276 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_247
timestamp 1666464484
transform 1 0 23828 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_253
timestamp 1666464484
transform 1 0 24380 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_256
timestamp 1666464484
transform 1 0 24656 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_262
timestamp 1666464484
transform 1 0 25208 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_268
timestamp 1666464484
transform 1 0 25760 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_271
timestamp 1666464484
transform 1 0 26036 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_277
timestamp 1666464484
transform 1 0 26588 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_283
timestamp 1666464484
transform 1 0 27140 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_286
timestamp 1666464484
transform 1 0 27416 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_292
timestamp 1666464484
transform 1 0 27968 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_298
timestamp 1666464484
transform 1 0 28520 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_301
timestamp 1666464484
transform 1 0 28796 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_307
timestamp 1666464484
transform 1 0 29348 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_313
timestamp 1666464484
transform 1 0 29900 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_316
timestamp 1666464484
transform 1 0 30176 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_322
timestamp 1666464484
transform 1 0 30728 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_328
timestamp 1666464484
transform 1 0 31280 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_331
timestamp 1666464484
transform 1 0 31556 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_343
timestamp 1666464484
transform 1 0 32660 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_346
timestamp 1666464484
transform 1 0 32936 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_354
timestamp 1666464484
transform 1 0 33672 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_101_361
timestamp 1666464484
transform 1 0 34316 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_369
timestamp 1666464484
transform 1 0 35052 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_101_376
timestamp 1666464484
transform 1 0 35696 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_388
timestamp 1666464484
transform 1 0 36800 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_391
timestamp 1666464484
transform 1 0 37076 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_403
timestamp 1666464484
transform 1 0 38180 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_406
timestamp 1666464484
transform 1 0 38456 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_418
timestamp 1666464484
transform 1 0 39560 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_421
timestamp 1666464484
transform 1 0 39836 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_430
timestamp 1666464484
transform 1 0 40664 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_434
timestamp 1666464484
transform 1 0 41032 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_436
timestamp 1666464484
transform 1 0 41216 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_101_448
timestamp 1666464484
transform 1 0 42320 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_451
timestamp 1666464484
transform 1 0 42596 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_463
timestamp 1666464484
transform 1 0 43700 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_466
timestamp 1666464484
transform 1 0 43976 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_474
timestamp 1666464484
transform 1 0 44712 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_101_481
timestamp 1666464484
transform 1 0 45356 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_488
timestamp 1666464484
transform 1 0 46000 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_494
timestamp 1666464484
transform 1 0 46552 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_496
timestamp 1666464484
transform 1 0 46736 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_508
timestamp 1666464484
transform 1 0 47840 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_511
timestamp 1666464484
transform 1 0 48116 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_523
timestamp 1666464484
transform 1 0 49220 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_526
timestamp 1666464484
transform 1 0 49496 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_538
timestamp 1666464484
transform 1 0 50600 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_101_541
timestamp 1666464484
transform 1 0 50876 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_548
timestamp 1666464484
transform 1 0 51520 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_554
timestamp 1666464484
transform 1 0 52072 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_556
timestamp 1666464484
transform 1 0 52256 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_565
timestamp 1666464484
transform 1 0 53084 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_569
timestamp 1666464484
transform 1 0 53452 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_571
timestamp 1666464484
transform 1 0 53636 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_578
timestamp 1666464484
transform 1 0 54280 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_584
timestamp 1666464484
transform 1 0 54832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_586
timestamp 1666464484
transform 1 0 55016 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_593
timestamp 1666464484
transform 1 0 55660 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_599
timestamp 1666464484
transform 1 0 56212 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_601
timestamp 1666464484
transform 1 0 56396 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_606
timestamp 1666464484
transform 1 0 56856 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_614
timestamp 1666464484
transform 1 0 57592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_616
timestamp 1666464484
transform 1 0 57776 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_624
timestamp 1666464484
transform 1 0 58512 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666464484
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666464484
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666464484
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666464484
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666464484
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666464484
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666464484
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666464484
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666464484
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666464484
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666464484
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666464484
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666464484
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666464484
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666464484
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666464484
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666464484
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666464484
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666464484
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666464484
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666464484
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666464484
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666464484
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666464484
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666464484
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666464484
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666464484
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666464484
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666464484
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666464484
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666464484
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666464484
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666464484
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666464484
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666464484
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666464484
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1666464484
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1666464484
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1666464484
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1666464484
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1666464484
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1666464484
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1666464484
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1666464484
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1666464484
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1666464484
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1666464484
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1666464484
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1666464484
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1666464484
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1666464484
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1666464484
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1666464484
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1666464484
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1666464484
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1666464484
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1666464484
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1666464484
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1666464484
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1666464484
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1666464484
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1666464484
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1666464484
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1666464484
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1666464484
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1666464484
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1666464484
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1666464484
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1666464484
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1666464484
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1666464484
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1666464484
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1666464484
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1666464484
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 3864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 5244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 6624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 8004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 9384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 10764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 12144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 13524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 14904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 17664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 20424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 23184 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 24564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 25944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 27324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 28704 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 30084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 31464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 34224 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 35604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 36984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 38364 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 41124 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 42504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 43884 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 45264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 46644 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 48024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 49404 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 50784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 52164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 53544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 54924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 56304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 3864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 6624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 9384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 12144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 14904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 17664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 20424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 23184 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 25944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 28704 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 31464 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 34224 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 36984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 39744 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 42504 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 45264 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 48024 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 50784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 53544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 56304 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 5244 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 8004 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 13524 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 21804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 24564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 27324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 30084 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 32844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 35604 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 38364 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 41124 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 43884 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 46644 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 49404 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 52164 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 54924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 57684 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 3864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 6624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 9384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 12144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 14904 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 17664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 20424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 23184 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 25944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 28704 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 31464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 34224 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 36984 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 39744 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 42504 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 45264 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 48024 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 50784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 53544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 56304 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 5244 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 8004 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 10764 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 13524 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 21804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 24564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 27324 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 30084 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 32844 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 35604 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 38364 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 41124 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 43884 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 46644 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 49404 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 52164 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 54924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 57684 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 3864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 6624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 9384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 12144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 14904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 17664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 20424 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 23184 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 25944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 28704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 31464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 34224 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 36984 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 39744 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 42504 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 45264 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 48024 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 50784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 53544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 56304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 5244 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 8004 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 10764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 13524 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 21804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 24564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 27324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 30084 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 32844 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 35604 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 38364 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 41124 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 43884 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 46644 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 49404 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 52164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 54924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 57684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 3864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 6624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 9384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 12144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 14904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 17664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 20424 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 23184 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 25944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 28704 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 31464 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 34224 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 36984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 39744 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 42504 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 45264 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 48024 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 50784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 53544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 56304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 5244 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 8004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 10764 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 13524 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 21804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 24564 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 27324 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 30084 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 32844 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 35604 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 38364 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 41124 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 43884 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 46644 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 49404 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 52164 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 54924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 57684 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 3864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 6624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 9384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 12144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 14904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 17664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 20424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 23184 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 25944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 28704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 31464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 34224 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 36984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 42504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 45264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 48024 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 50784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 53544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 56304 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 5244 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 8004 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 10764 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 13524 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 21804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 24564 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 27324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 30084 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 32844 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 35604 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 38364 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 41124 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 43884 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 46644 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 49404 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 52164 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 54924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 57684 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 3864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 6624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 9384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 12144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 14904 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 17664 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 20424 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 23184 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 25944 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 28704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 31464 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 34224 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 36984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 42504 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 45264 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 48024 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 50784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 53544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 56304 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 5244 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 8004 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 10764 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 13524 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 21804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 24564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 27324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 30084 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 32844 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 35604 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 38364 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 41124 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 43884 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 46644 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 49404 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 52164 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 54924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 57684 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 3864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 6624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 9384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 12144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 14904 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 17664 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 20424 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 23184 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 25944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 28704 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 31464 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 34224 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 36984 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 39744 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 42504 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 45264 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 48024 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 50784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 53544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 56304 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 5244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 8004 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 10764 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 13524 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 21804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 24564 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 27324 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 30084 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 32844 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 35604 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 38364 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 41124 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 43884 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 46644 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 49404 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 52164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 54924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 57684 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 3864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 6624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 9384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 12144 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 14904 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 17664 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 20424 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 23184 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 25944 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 28704 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 31464 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 34224 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 36984 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 39744 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 42504 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 45264 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 48024 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 50784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 53544 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 56304 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 5244 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 8004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 10764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 13524 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 21804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 24564 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 27324 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 30084 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 32844 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666464484
transform 1 0 35604 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666464484
transform 1 0 38364 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666464484
transform 1 0 41124 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666464484
transform 1 0 43884 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666464484
transform 1 0 46644 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666464484
transform 1 0 49404 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666464484
transform 1 0 52164 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666464484
transform 1 0 54924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666464484
transform 1 0 57684 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666464484
transform 1 0 3864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666464484
transform 1 0 6624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666464484
transform 1 0 9384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666464484
transform 1 0 12144 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666464484
transform 1 0 14904 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666464484
transform 1 0 17664 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666464484
transform 1 0 20424 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666464484
transform 1 0 23184 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666464484
transform 1 0 25944 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666464484
transform 1 0 28704 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666464484
transform 1 0 31464 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666464484
transform 1 0 34224 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666464484
transform 1 0 36984 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666464484
transform 1 0 39744 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666464484
transform 1 0 42504 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666464484
transform 1 0 45264 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666464484
transform 1 0 48024 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666464484
transform 1 0 50784 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666464484
transform 1 0 53544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666464484
transform 1 0 56304 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666464484
transform 1 0 5244 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666464484
transform 1 0 8004 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666464484
transform 1 0 10764 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666464484
transform 1 0 13524 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666464484
transform 1 0 21804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666464484
transform 1 0 24564 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666464484
transform 1 0 27324 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666464484
transform 1 0 30084 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666464484
transform 1 0 32844 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666464484
transform 1 0 35604 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666464484
transform 1 0 38364 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666464484
transform 1 0 41124 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666464484
transform 1 0 43884 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666464484
transform 1 0 46644 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666464484
transform 1 0 49404 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666464484
transform 1 0 52164 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666464484
transform 1 0 54924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666464484
transform 1 0 57684 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666464484
transform 1 0 3864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666464484
transform 1 0 6624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666464484
transform 1 0 9384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666464484
transform 1 0 12144 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666464484
transform 1 0 14904 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666464484
transform 1 0 17664 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666464484
transform 1 0 20424 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666464484
transform 1 0 23184 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666464484
transform 1 0 25944 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666464484
transform 1 0 28704 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666464484
transform 1 0 31464 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666464484
transform 1 0 34224 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666464484
transform 1 0 36984 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666464484
transform 1 0 39744 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666464484
transform 1 0 42504 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666464484
transform 1 0 45264 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666464484
transform 1 0 48024 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666464484
transform 1 0 50784 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666464484
transform 1 0 53544 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666464484
transform 1 0 56304 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666464484
transform 1 0 2484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666464484
transform 1 0 5244 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666464484
transform 1 0 8004 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666464484
transform 1 0 10764 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666464484
transform 1 0 13524 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666464484
transform 1 0 21804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666464484
transform 1 0 24564 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666464484
transform 1 0 27324 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666464484
transform 1 0 30084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666464484
transform 1 0 32844 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666464484
transform 1 0 35604 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666464484
transform 1 0 38364 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666464484
transform 1 0 41124 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666464484
transform 1 0 43884 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666464484
transform 1 0 46644 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666464484
transform 1 0 49404 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666464484
transform 1 0 52164 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666464484
transform 1 0 54924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666464484
transform 1 0 57684 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666464484
transform 1 0 3864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666464484
transform 1 0 6624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666464484
transform 1 0 9384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666464484
transform 1 0 12144 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666464484
transform 1 0 14904 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666464484
transform 1 0 17664 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666464484
transform 1 0 20424 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666464484
transform 1 0 23184 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666464484
transform 1 0 25944 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666464484
transform 1 0 28704 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666464484
transform 1 0 31464 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666464484
transform 1 0 34224 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666464484
transform 1 0 36984 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666464484
transform 1 0 39744 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666464484
transform 1 0 42504 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666464484
transform 1 0 45264 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666464484
transform 1 0 48024 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666464484
transform 1 0 50784 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666464484
transform 1 0 53544 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666464484
transform 1 0 56304 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666464484
transform 1 0 2484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666464484
transform 1 0 5244 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666464484
transform 1 0 8004 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666464484
transform 1 0 10764 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666464484
transform 1 0 13524 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666464484
transform 1 0 21804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666464484
transform 1 0 24564 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666464484
transform 1 0 27324 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666464484
transform 1 0 30084 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666464484
transform 1 0 32844 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666464484
transform 1 0 35604 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666464484
transform 1 0 38364 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666464484
transform 1 0 41124 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666464484
transform 1 0 43884 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666464484
transform 1 0 46644 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666464484
transform 1 0 49404 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666464484
transform 1 0 52164 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666464484
transform 1 0 54924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666464484
transform 1 0 57684 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666464484
transform 1 0 3864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666464484
transform 1 0 6624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666464484
transform 1 0 9384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666464484
transform 1 0 12144 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666464484
transform 1 0 14904 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666464484
transform 1 0 17664 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666464484
transform 1 0 20424 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666464484
transform 1 0 23184 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666464484
transform 1 0 25944 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666464484
transform 1 0 28704 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666464484
transform 1 0 31464 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666464484
transform 1 0 34224 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666464484
transform 1 0 36984 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666464484
transform 1 0 39744 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666464484
transform 1 0 42504 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666464484
transform 1 0 45264 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666464484
transform 1 0 48024 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666464484
transform 1 0 50784 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666464484
transform 1 0 53544 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666464484
transform 1 0 56304 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666464484
transform 1 0 5244 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666464484
transform 1 0 8004 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666464484
transform 1 0 10764 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666464484
transform 1 0 13524 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666464484
transform 1 0 21804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666464484
transform 1 0 24564 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666464484
transform 1 0 27324 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666464484
transform 1 0 30084 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666464484
transform 1 0 32844 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666464484
transform 1 0 35604 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666464484
transform 1 0 38364 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666464484
transform 1 0 41124 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666464484
transform 1 0 43884 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666464484
transform 1 0 46644 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666464484
transform 1 0 49404 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666464484
transform 1 0 52164 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666464484
transform 1 0 54924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666464484
transform 1 0 57684 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666464484
transform 1 0 3864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666464484
transform 1 0 6624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666464484
transform 1 0 9384 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666464484
transform 1 0 12144 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666464484
transform 1 0 14904 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666464484
transform 1 0 17664 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666464484
transform 1 0 20424 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666464484
transform 1 0 23184 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666464484
transform 1 0 25944 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666464484
transform 1 0 28704 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666464484
transform 1 0 31464 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666464484
transform 1 0 34224 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666464484
transform 1 0 36984 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666464484
transform 1 0 39744 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666464484
transform 1 0 42504 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666464484
transform 1 0 45264 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666464484
transform 1 0 48024 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666464484
transform 1 0 50784 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666464484
transform 1 0 53544 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666464484
transform 1 0 56304 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666464484
transform 1 0 5244 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666464484
transform 1 0 8004 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666464484
transform 1 0 10764 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666464484
transform 1 0 13524 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666464484
transform 1 0 21804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666464484
transform 1 0 24564 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666464484
transform 1 0 27324 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666464484
transform 1 0 30084 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666464484
transform 1 0 32844 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666464484
transform 1 0 35604 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666464484
transform 1 0 38364 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666464484
transform 1 0 41124 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666464484
transform 1 0 43884 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666464484
transform 1 0 46644 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666464484
transform 1 0 49404 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666464484
transform 1 0 52164 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666464484
transform 1 0 54924 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666464484
transform 1 0 57684 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666464484
transform 1 0 3864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666464484
transform 1 0 6624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666464484
transform 1 0 9384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666464484
transform 1 0 12144 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666464484
transform 1 0 14904 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666464484
transform 1 0 17664 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666464484
transform 1 0 20424 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666464484
transform 1 0 23184 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666464484
transform 1 0 25944 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666464484
transform 1 0 28704 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666464484
transform 1 0 31464 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666464484
transform 1 0 34224 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666464484
transform 1 0 36984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666464484
transform 1 0 39744 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666464484
transform 1 0 42504 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666464484
transform 1 0 45264 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666464484
transform 1 0 48024 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666464484
transform 1 0 50784 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666464484
transform 1 0 53544 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666464484
transform 1 0 56304 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666464484
transform 1 0 2484 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666464484
transform 1 0 5244 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666464484
transform 1 0 8004 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666464484
transform 1 0 10764 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666464484
transform 1 0 13524 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666464484
transform 1 0 21804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666464484
transform 1 0 24564 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666464484
transform 1 0 27324 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666464484
transform 1 0 30084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666464484
transform 1 0 32844 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666464484
transform 1 0 35604 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666464484
transform 1 0 38364 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666464484
transform 1 0 41124 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666464484
transform 1 0 43884 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666464484
transform 1 0 46644 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666464484
transform 1 0 49404 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666464484
transform 1 0 52164 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666464484
transform 1 0 54924 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666464484
transform 1 0 57684 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666464484
transform 1 0 3864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666464484
transform 1 0 6624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666464484
transform 1 0 9384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666464484
transform 1 0 12144 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666464484
transform 1 0 14904 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666464484
transform 1 0 17664 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666464484
transform 1 0 20424 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666464484
transform 1 0 23184 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666464484
transform 1 0 25944 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666464484
transform 1 0 28704 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666464484
transform 1 0 31464 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666464484
transform 1 0 34224 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666464484
transform 1 0 36984 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666464484
transform 1 0 39744 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666464484
transform 1 0 42504 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666464484
transform 1 0 45264 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666464484
transform 1 0 48024 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666464484
transform 1 0 50784 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666464484
transform 1 0 53544 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666464484
transform 1 0 56304 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666464484
transform 1 0 5244 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666464484
transform 1 0 8004 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666464484
transform 1 0 10764 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666464484
transform 1 0 13524 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666464484
transform 1 0 21804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666464484
transform 1 0 24564 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666464484
transform 1 0 27324 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666464484
transform 1 0 30084 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666464484
transform 1 0 32844 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666464484
transform 1 0 35604 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666464484
transform 1 0 38364 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666464484
transform 1 0 41124 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666464484
transform 1 0 43884 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666464484
transform 1 0 46644 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666464484
transform 1 0 49404 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666464484
transform 1 0 52164 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666464484
transform 1 0 54924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666464484
transform 1 0 57684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666464484
transform 1 0 3864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666464484
transform 1 0 6624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666464484
transform 1 0 9384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666464484
transform 1 0 12144 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666464484
transform 1 0 14904 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666464484
transform 1 0 17664 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666464484
transform 1 0 20424 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666464484
transform 1 0 23184 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666464484
transform 1 0 25944 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666464484
transform 1 0 28704 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666464484
transform 1 0 31464 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666464484
transform 1 0 34224 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666464484
transform 1 0 36984 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666464484
transform 1 0 39744 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666464484
transform 1 0 42504 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666464484
transform 1 0 45264 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666464484
transform 1 0 48024 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666464484
transform 1 0 50784 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666464484
transform 1 0 53544 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666464484
transform 1 0 56304 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666464484
transform 1 0 5244 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666464484
transform 1 0 8004 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666464484
transform 1 0 10764 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666464484
transform 1 0 13524 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666464484
transform 1 0 21804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666464484
transform 1 0 24564 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666464484
transform 1 0 27324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666464484
transform 1 0 30084 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666464484
transform 1 0 32844 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666464484
transform 1 0 35604 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666464484
transform 1 0 38364 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666464484
transform 1 0 41124 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666464484
transform 1 0 43884 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666464484
transform 1 0 46644 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666464484
transform 1 0 49404 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666464484
transform 1 0 52164 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666464484
transform 1 0 54924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666464484
transform 1 0 57684 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666464484
transform 1 0 3864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666464484
transform 1 0 6624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666464484
transform 1 0 9384 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666464484
transform 1 0 12144 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666464484
transform 1 0 14904 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666464484
transform 1 0 17664 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666464484
transform 1 0 20424 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666464484
transform 1 0 23184 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666464484
transform 1 0 25944 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666464484
transform 1 0 28704 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666464484
transform 1 0 31464 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666464484
transform 1 0 34224 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666464484
transform 1 0 36984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666464484
transform 1 0 39744 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666464484
transform 1 0 42504 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666464484
transform 1 0 45264 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666464484
transform 1 0 48024 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666464484
transform 1 0 50784 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666464484
transform 1 0 53544 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666464484
transform 1 0 56304 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666464484
transform 1 0 5244 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666464484
transform 1 0 8004 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666464484
transform 1 0 10764 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666464484
transform 1 0 13524 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666464484
transform 1 0 21804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666464484
transform 1 0 24564 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666464484
transform 1 0 27324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1666464484
transform 1 0 30084 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1666464484
transform 1 0 32844 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1666464484
transform 1 0 35604 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1666464484
transform 1 0 38364 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1666464484
transform 1 0 41124 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1666464484
transform 1 0 43884 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1666464484
transform 1 0 46644 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1666464484
transform 1 0 49404 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1666464484
transform 1 0 52164 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1666464484
transform 1 0 54924 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1666464484
transform 1 0 57684 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1666464484
transform 1 0 3864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1666464484
transform 1 0 6624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1666464484
transform 1 0 9384 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1666464484
transform 1 0 12144 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1666464484
transform 1 0 14904 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1666464484
transform 1 0 17664 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1666464484
transform 1 0 20424 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1666464484
transform 1 0 23184 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1666464484
transform 1 0 25944 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1666464484
transform 1 0 28704 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1666464484
transform 1 0 31464 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1666464484
transform 1 0 34224 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1666464484
transform 1 0 36984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1666464484
transform 1 0 39744 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1666464484
transform 1 0 42504 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1666464484
transform 1 0 45264 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1666464484
transform 1 0 48024 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1666464484
transform 1 0 50784 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1666464484
transform 1 0 53544 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1666464484
transform 1 0 56304 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1666464484
transform 1 0 5244 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1666464484
transform 1 0 8004 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1666464484
transform 1 0 10764 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1666464484
transform 1 0 13524 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1666464484
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1666464484
transform 1 0 21804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1666464484
transform 1 0 24564 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1666464484
transform 1 0 27324 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1666464484
transform 1 0 30084 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1666464484
transform 1 0 32844 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1666464484
transform 1 0 35604 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1666464484
transform 1 0 38364 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1666464484
transform 1 0 41124 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1666464484
transform 1 0 43884 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1666464484
transform 1 0 46644 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1666464484
transform 1 0 49404 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1666464484
transform 1 0 52164 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1666464484
transform 1 0 54924 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1666464484
transform 1 0 57684 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1666464484
transform 1 0 3864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1666464484
transform 1 0 6624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1666464484
transform 1 0 9384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1666464484
transform 1 0 12144 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1666464484
transform 1 0 14904 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1666464484
transform 1 0 17664 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1666464484
transform 1 0 20424 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1666464484
transform 1 0 23184 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1666464484
transform 1 0 25944 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1666464484
transform 1 0 28704 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1666464484
transform 1 0 31464 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1666464484
transform 1 0 34224 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1666464484
transform 1 0 36984 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1666464484
transform 1 0 39744 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1666464484
transform 1 0 42504 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1666464484
transform 1 0 45264 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1666464484
transform 1 0 48024 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1666464484
transform 1 0 50784 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1666464484
transform 1 0 53544 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1666464484
transform 1 0 56304 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1666464484
transform 1 0 5244 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1666464484
transform 1 0 8004 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1666464484
transform 1 0 10764 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1666464484
transform 1 0 13524 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1666464484
transform 1 0 16284 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1666464484
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1666464484
transform 1 0 21804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1666464484
transform 1 0 24564 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1666464484
transform 1 0 27324 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1666464484
transform 1 0 30084 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1666464484
transform 1 0 32844 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1666464484
transform 1 0 35604 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1666464484
transform 1 0 38364 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1666464484
transform 1 0 41124 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1666464484
transform 1 0 43884 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1666464484
transform 1 0 46644 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1666464484
transform 1 0 49404 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1666464484
transform 1 0 52164 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1666464484
transform 1 0 54924 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1666464484
transform 1 0 57684 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1666464484
transform 1 0 3864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1666464484
transform 1 0 6624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1666464484
transform 1 0 9384 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1666464484
transform 1 0 12144 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1666464484
transform 1 0 14904 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1666464484
transform 1 0 17664 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1666464484
transform 1 0 20424 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1666464484
transform 1 0 23184 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1666464484
transform 1 0 25944 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1666464484
transform 1 0 28704 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1666464484
transform 1 0 31464 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1666464484
transform 1 0 34224 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1666464484
transform 1 0 36984 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1666464484
transform 1 0 39744 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1666464484
transform 1 0 42504 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1666464484
transform 1 0 45264 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1666464484
transform 1 0 48024 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1666464484
transform 1 0 50784 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1666464484
transform 1 0 53544 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1666464484
transform 1 0 56304 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1666464484
transform 1 0 2484 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1666464484
transform 1 0 5244 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1666464484
transform 1 0 8004 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1666464484
transform 1 0 10764 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1666464484
transform 1 0 13524 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1666464484
transform 1 0 16284 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1666464484
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1666464484
transform 1 0 21804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1666464484
transform 1 0 24564 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1666464484
transform 1 0 27324 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1666464484
transform 1 0 30084 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1666464484
transform 1 0 32844 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1666464484
transform 1 0 35604 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1666464484
transform 1 0 38364 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1666464484
transform 1 0 41124 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1666464484
transform 1 0 43884 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1666464484
transform 1 0 46644 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1666464484
transform 1 0 49404 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1666464484
transform 1 0 52164 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1666464484
transform 1 0 54924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1666464484
transform 1 0 57684 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1666464484
transform 1 0 3864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1666464484
transform 1 0 6624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1666464484
transform 1 0 9384 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1666464484
transform 1 0 12144 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1666464484
transform 1 0 14904 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1666464484
transform 1 0 17664 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1666464484
transform 1 0 20424 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1666464484
transform 1 0 23184 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1666464484
transform 1 0 25944 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1666464484
transform 1 0 28704 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1666464484
transform 1 0 31464 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1666464484
transform 1 0 34224 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1666464484
transform 1 0 36984 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1666464484
transform 1 0 39744 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1666464484
transform 1 0 42504 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1666464484
transform 1 0 45264 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1666464484
transform 1 0 48024 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1666464484
transform 1 0 50784 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1666464484
transform 1 0 53544 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1666464484
transform 1 0 56304 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1666464484
transform 1 0 5244 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1666464484
transform 1 0 8004 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1666464484
transform 1 0 10764 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1666464484
transform 1 0 13524 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1666464484
transform 1 0 16284 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1666464484
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1666464484
transform 1 0 21804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1666464484
transform 1 0 24564 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1666464484
transform 1 0 27324 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1666464484
transform 1 0 30084 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1666464484
transform 1 0 32844 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1666464484
transform 1 0 35604 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1666464484
transform 1 0 38364 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1666464484
transform 1 0 41124 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1666464484
transform 1 0 43884 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1666464484
transform 1 0 46644 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1666464484
transform 1 0 49404 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1666464484
transform 1 0 52164 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1666464484
transform 1 0 54924 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1666464484
transform 1 0 57684 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1666464484
transform 1 0 3864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1666464484
transform 1 0 6624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1666464484
transform 1 0 9384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1666464484
transform 1 0 12144 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1666464484
transform 1 0 14904 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1666464484
transform 1 0 17664 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1666464484
transform 1 0 20424 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1666464484
transform 1 0 23184 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1666464484
transform 1 0 25944 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1666464484
transform 1 0 28704 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1666464484
transform 1 0 31464 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1666464484
transform 1 0 34224 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1666464484
transform 1 0 36984 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1666464484
transform 1 0 39744 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1666464484
transform 1 0 42504 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1666464484
transform 1 0 45264 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1666464484
transform 1 0 48024 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1666464484
transform 1 0 50784 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1666464484
transform 1 0 53544 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1666464484
transform 1 0 56304 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1666464484
transform 1 0 5244 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1666464484
transform 1 0 8004 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1666464484
transform 1 0 10764 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1666464484
transform 1 0 13524 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1666464484
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1666464484
transform 1 0 21804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1666464484
transform 1 0 24564 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1666464484
transform 1 0 27324 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1666464484
transform 1 0 30084 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1666464484
transform 1 0 32844 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1666464484
transform 1 0 35604 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1666464484
transform 1 0 38364 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1666464484
transform 1 0 41124 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1666464484
transform 1 0 43884 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1666464484
transform 1 0 46644 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1666464484
transform 1 0 49404 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1666464484
transform 1 0 52164 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1666464484
transform 1 0 54924 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1666464484
transform 1 0 57684 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1666464484
transform 1 0 3864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1666464484
transform 1 0 6624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1666464484
transform 1 0 9384 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1666464484
transform 1 0 12144 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1666464484
transform 1 0 14904 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1666464484
transform 1 0 17664 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1666464484
transform 1 0 20424 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1666464484
transform 1 0 23184 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1666464484
transform 1 0 25944 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1666464484
transform 1 0 28704 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1666464484
transform 1 0 31464 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1666464484
transform 1 0 34224 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1666464484
transform 1 0 36984 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1666464484
transform 1 0 39744 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1666464484
transform 1 0 42504 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1666464484
transform 1 0 45264 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1666464484
transform 1 0 48024 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1666464484
transform 1 0 50784 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1666464484
transform 1 0 53544 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1666464484
transform 1 0 56304 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1666464484
transform 1 0 5244 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1666464484
transform 1 0 8004 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1666464484
transform 1 0 10764 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1666464484
transform 1 0 13524 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1666464484
transform 1 0 16284 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1666464484
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1666464484
transform 1 0 21804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1666464484
transform 1 0 24564 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1666464484
transform 1 0 27324 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1666464484
transform 1 0 30084 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1666464484
transform 1 0 32844 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1666464484
transform 1 0 35604 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1666464484
transform 1 0 38364 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1666464484
transform 1 0 41124 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1666464484
transform 1 0 43884 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1666464484
transform 1 0 46644 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1666464484
transform 1 0 49404 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1666464484
transform 1 0 52164 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1666464484
transform 1 0 54924 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1666464484
transform 1 0 57684 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1666464484
transform 1 0 3864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1666464484
transform 1 0 6624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1666464484
transform 1 0 9384 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1666464484
transform 1 0 12144 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1666464484
transform 1 0 14904 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1666464484
transform 1 0 17664 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1666464484
transform 1 0 20424 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1666464484
transform 1 0 23184 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1666464484
transform 1 0 25944 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1666464484
transform 1 0 28704 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1666464484
transform 1 0 31464 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1666464484
transform 1 0 34224 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1666464484
transform 1 0 36984 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1666464484
transform 1 0 39744 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1666464484
transform 1 0 42504 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1666464484
transform 1 0 45264 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1666464484
transform 1 0 48024 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1666464484
transform 1 0 50784 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1666464484
transform 1 0 53544 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1666464484
transform 1 0 56304 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1666464484
transform 1 0 5244 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1666464484
transform 1 0 8004 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1666464484
transform 1 0 10764 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1666464484
transform 1 0 13524 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1666464484
transform 1 0 16284 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1666464484
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1666464484
transform 1 0 21804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1666464484
transform 1 0 24564 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1666464484
transform 1 0 27324 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1666464484
transform 1 0 30084 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1666464484
transform 1 0 32844 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1666464484
transform 1 0 35604 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1666464484
transform 1 0 38364 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1666464484
transform 1 0 41124 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1666464484
transform 1 0 43884 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1666464484
transform 1 0 46644 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1666464484
transform 1 0 49404 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1666464484
transform 1 0 52164 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1666464484
transform 1 0 54924 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1666464484
transform 1 0 57684 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1666464484
transform 1 0 3864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1666464484
transform 1 0 6624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1666464484
transform 1 0 9384 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1666464484
transform 1 0 12144 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1666464484
transform 1 0 14904 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1666464484
transform 1 0 17664 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1666464484
transform 1 0 20424 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1666464484
transform 1 0 23184 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1666464484
transform 1 0 25944 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1666464484
transform 1 0 28704 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1666464484
transform 1 0 31464 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1666464484
transform 1 0 34224 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1666464484
transform 1 0 36984 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1666464484
transform 1 0 39744 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1666464484
transform 1 0 42504 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1666464484
transform 1 0 45264 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1666464484
transform 1 0 48024 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1666464484
transform 1 0 50784 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1666464484
transform 1 0 53544 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1666464484
transform 1 0 56304 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1666464484
transform 1 0 5244 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1666464484
transform 1 0 8004 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1666464484
transform 1 0 10764 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1666464484
transform 1 0 13524 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1666464484
transform 1 0 16284 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1666464484
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1666464484
transform 1 0 21804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1666464484
transform 1 0 24564 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1666464484
transform 1 0 27324 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1666464484
transform 1 0 30084 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1666464484
transform 1 0 32844 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1666464484
transform 1 0 35604 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1666464484
transform 1 0 38364 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1666464484
transform 1 0 41124 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1666464484
transform 1 0 43884 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1666464484
transform 1 0 46644 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1666464484
transform 1 0 49404 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1666464484
transform 1 0 52164 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1666464484
transform 1 0 54924 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1666464484
transform 1 0 57684 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1666464484
transform 1 0 3864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1666464484
transform 1 0 6624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1666464484
transform 1 0 9384 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1666464484
transform 1 0 12144 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1666464484
transform 1 0 14904 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1666464484
transform 1 0 17664 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1666464484
transform 1 0 20424 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1666464484
transform 1 0 23184 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1666464484
transform 1 0 25944 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1666464484
transform 1 0 28704 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1666464484
transform 1 0 31464 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1666464484
transform 1 0 34224 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1666464484
transform 1 0 36984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1666464484
transform 1 0 39744 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1666464484
transform 1 0 42504 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1666464484
transform 1 0 45264 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1666464484
transform 1 0 48024 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1666464484
transform 1 0 50784 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1666464484
transform 1 0 53544 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1666464484
transform 1 0 56304 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1666464484
transform 1 0 5244 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1666464484
transform 1 0 8004 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1666464484
transform 1 0 10764 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1666464484
transform 1 0 13524 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1666464484
transform 1 0 16284 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1666464484
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1666464484
transform 1 0 21804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1666464484
transform 1 0 24564 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1666464484
transform 1 0 27324 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1666464484
transform 1 0 30084 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1666464484
transform 1 0 32844 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1666464484
transform 1 0 35604 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1666464484
transform 1 0 38364 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1666464484
transform 1 0 41124 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1666464484
transform 1 0 43884 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1666464484
transform 1 0 46644 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1666464484
transform 1 0 49404 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1666464484
transform 1 0 52164 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1666464484
transform 1 0 54924 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1666464484
transform 1 0 57684 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1666464484
transform 1 0 3864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1666464484
transform 1 0 6624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1666464484
transform 1 0 9384 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1666464484
transform 1 0 12144 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1666464484
transform 1 0 14904 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1666464484
transform 1 0 17664 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1666464484
transform 1 0 20424 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1666464484
transform 1 0 23184 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1666464484
transform 1 0 25944 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1666464484
transform 1 0 28704 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1666464484
transform 1 0 31464 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1666464484
transform 1 0 34224 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1666464484
transform 1 0 36984 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1666464484
transform 1 0 39744 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1666464484
transform 1 0 42504 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1666464484
transform 1 0 45264 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1666464484
transform 1 0 48024 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1666464484
transform 1 0 50784 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1666464484
transform 1 0 53544 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1666464484
transform 1 0 56304 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1666464484
transform 1 0 2484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1666464484
transform 1 0 5244 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1666464484
transform 1 0 8004 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1666464484
transform 1 0 10764 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1666464484
transform 1 0 13524 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1666464484
transform 1 0 16284 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1666464484
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1666464484
transform 1 0 21804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1666464484
transform 1 0 24564 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1666464484
transform 1 0 27324 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1666464484
transform 1 0 30084 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1666464484
transform 1 0 32844 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1666464484
transform 1 0 35604 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1666464484
transform 1 0 38364 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1666464484
transform 1 0 41124 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1666464484
transform 1 0 43884 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1666464484
transform 1 0 46644 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1666464484
transform 1 0 49404 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1666464484
transform 1 0 52164 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1666464484
transform 1 0 54924 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1666464484
transform 1 0 57684 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1666464484
transform 1 0 3864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1666464484
transform 1 0 6624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1666464484
transform 1 0 9384 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1666464484
transform 1 0 12144 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1666464484
transform 1 0 14904 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1666464484
transform 1 0 17664 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1666464484
transform 1 0 20424 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1666464484
transform 1 0 23184 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1666464484
transform 1 0 25944 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1666464484
transform 1 0 28704 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1666464484
transform 1 0 31464 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1666464484
transform 1 0 34224 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1666464484
transform 1 0 36984 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1666464484
transform 1 0 39744 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1666464484
transform 1 0 42504 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1666464484
transform 1 0 45264 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1666464484
transform 1 0 48024 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1666464484
transform 1 0 50784 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1666464484
transform 1 0 53544 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1666464484
transform 1 0 56304 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1666464484
transform 1 0 2484 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1666464484
transform 1 0 5244 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1666464484
transform 1 0 8004 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1666464484
transform 1 0 10764 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1666464484
transform 1 0 13524 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1666464484
transform 1 0 16284 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1666464484
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1666464484
transform 1 0 21804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1666464484
transform 1 0 24564 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1666464484
transform 1 0 27324 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1666464484
transform 1 0 30084 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1666464484
transform 1 0 32844 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1666464484
transform 1 0 35604 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1666464484
transform 1 0 38364 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1666464484
transform 1 0 41124 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1666464484
transform 1 0 43884 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1666464484
transform 1 0 46644 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1666464484
transform 1 0 49404 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1666464484
transform 1 0 52164 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1666464484
transform 1 0 54924 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1666464484
transform 1 0 57684 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1666464484
transform 1 0 3864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1666464484
transform 1 0 6624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1666464484
transform 1 0 9384 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1666464484
transform 1 0 12144 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1666464484
transform 1 0 14904 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1666464484
transform 1 0 17664 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1666464484
transform 1 0 20424 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1666464484
transform 1 0 23184 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1666464484
transform 1 0 25944 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1666464484
transform 1 0 28704 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1666464484
transform 1 0 31464 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1666464484
transform 1 0 34224 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1666464484
transform 1 0 36984 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1666464484
transform 1 0 39744 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1666464484
transform 1 0 42504 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1666464484
transform 1 0 45264 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1666464484
transform 1 0 48024 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1666464484
transform 1 0 50784 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1666464484
transform 1 0 53544 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1666464484
transform 1 0 56304 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1666464484
transform 1 0 2484 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1666464484
transform 1 0 5244 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1666464484
transform 1 0 8004 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1666464484
transform 1 0 10764 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1666464484
transform 1 0 13524 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1666464484
transform 1 0 16284 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1666464484
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1666464484
transform 1 0 21804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1666464484
transform 1 0 24564 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1666464484
transform 1 0 27324 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1666464484
transform 1 0 30084 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1666464484
transform 1 0 32844 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1666464484
transform 1 0 35604 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1666464484
transform 1 0 38364 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1666464484
transform 1 0 41124 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1666464484
transform 1 0 43884 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1666464484
transform 1 0 46644 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1666464484
transform 1 0 49404 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1666464484
transform 1 0 52164 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1666464484
transform 1 0 54924 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1666464484
transform 1 0 57684 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1666464484
transform 1 0 3864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1666464484
transform 1 0 6624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1666464484
transform 1 0 9384 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1666464484
transform 1 0 12144 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1666464484
transform 1 0 14904 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1666464484
transform 1 0 17664 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1666464484
transform 1 0 20424 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1666464484
transform 1 0 23184 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1666464484
transform 1 0 25944 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1666464484
transform 1 0 28704 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1666464484
transform 1 0 31464 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1666464484
transform 1 0 34224 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1666464484
transform 1 0 36984 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1666464484
transform 1 0 39744 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1666464484
transform 1 0 42504 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1666464484
transform 1 0 45264 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1666464484
transform 1 0 48024 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1666464484
transform 1 0 50784 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1666464484
transform 1 0 53544 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1666464484
transform 1 0 56304 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1666464484
transform 1 0 2484 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1666464484
transform 1 0 5244 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1666464484
transform 1 0 8004 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1666464484
transform 1 0 10764 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1666464484
transform 1 0 13524 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1666464484
transform 1 0 16284 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1666464484
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1666464484
transform 1 0 21804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1666464484
transform 1 0 24564 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1666464484
transform 1 0 27324 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1666464484
transform 1 0 30084 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1666464484
transform 1 0 32844 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1666464484
transform 1 0 35604 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1666464484
transform 1 0 38364 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1666464484
transform 1 0 41124 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1666464484
transform 1 0 43884 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1666464484
transform 1 0 46644 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1666464484
transform 1 0 49404 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1666464484
transform 1 0 52164 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1666464484
transform 1 0 54924 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1666464484
transform 1 0 57684 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1666464484
transform 1 0 3864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1666464484
transform 1 0 6624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1666464484
transform 1 0 9384 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1666464484
transform 1 0 12144 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1666464484
transform 1 0 14904 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1666464484
transform 1 0 17664 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1666464484
transform 1 0 20424 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1666464484
transform 1 0 23184 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1666464484
transform 1 0 25944 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1666464484
transform 1 0 28704 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1666464484
transform 1 0 31464 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1666464484
transform 1 0 34224 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1666464484
transform 1 0 36984 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1666464484
transform 1 0 39744 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1666464484
transform 1 0 42504 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1666464484
transform 1 0 45264 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1666464484
transform 1 0 48024 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1666464484
transform 1 0 50784 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1666464484
transform 1 0 53544 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1666464484
transform 1 0 56304 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1666464484
transform 1 0 2484 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1666464484
transform 1 0 5244 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1666464484
transform 1 0 8004 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1666464484
transform 1 0 10764 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1666464484
transform 1 0 13524 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1666464484
transform 1 0 16284 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1666464484
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1666464484
transform 1 0 21804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1666464484
transform 1 0 24564 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1666464484
transform 1 0 27324 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1666464484
transform 1 0 30084 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1666464484
transform 1 0 32844 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1666464484
transform 1 0 35604 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1666464484
transform 1 0 38364 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1666464484
transform 1 0 41124 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1666464484
transform 1 0 43884 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1666464484
transform 1 0 46644 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1666464484
transform 1 0 49404 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1666464484
transform 1 0 52164 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1666464484
transform 1 0 54924 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1666464484
transform 1 0 57684 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1666464484
transform 1 0 3864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1666464484
transform 1 0 6624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1666464484
transform 1 0 9384 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1666464484
transform 1 0 12144 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1666464484
transform 1 0 14904 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1666464484
transform 1 0 17664 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1666464484
transform 1 0 20424 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1666464484
transform 1 0 23184 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1666464484
transform 1 0 25944 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1666464484
transform 1 0 28704 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1666464484
transform 1 0 31464 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1666464484
transform 1 0 34224 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1666464484
transform 1 0 36984 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1666464484
transform 1 0 39744 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1666464484
transform 1 0 42504 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1666464484
transform 1 0 45264 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1666464484
transform 1 0 48024 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1666464484
transform 1 0 50784 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1666464484
transform 1 0 53544 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1666464484
transform 1 0 56304 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1666464484
transform 1 0 2484 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1666464484
transform 1 0 5244 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1666464484
transform 1 0 8004 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1666464484
transform 1 0 10764 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1666464484
transform 1 0 13524 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1666464484
transform 1 0 16284 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1666464484
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1666464484
transform 1 0 21804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1666464484
transform 1 0 24564 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1666464484
transform 1 0 27324 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1666464484
transform 1 0 30084 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1666464484
transform 1 0 32844 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1666464484
transform 1 0 35604 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1666464484
transform 1 0 38364 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1666464484
transform 1 0 41124 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1666464484
transform 1 0 43884 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1666464484
transform 1 0 46644 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1666464484
transform 1 0 49404 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1666464484
transform 1 0 52164 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1666464484
transform 1 0 54924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1666464484
transform 1 0 57684 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1666464484
transform 1 0 3864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1666464484
transform 1 0 6624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1666464484
transform 1 0 9384 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1666464484
transform 1 0 12144 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1666464484
transform 1 0 14904 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1666464484
transform 1 0 17664 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1666464484
transform 1 0 20424 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1666464484
transform 1 0 23184 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1666464484
transform 1 0 25944 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1666464484
transform 1 0 28704 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1666464484
transform 1 0 31464 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1666464484
transform 1 0 34224 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1666464484
transform 1 0 36984 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1666464484
transform 1 0 39744 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1666464484
transform 1 0 42504 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1666464484
transform 1 0 45264 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1666464484
transform 1 0 48024 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1666464484
transform 1 0 50784 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1666464484
transform 1 0 53544 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1666464484
transform 1 0 56304 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1666464484
transform 1 0 2484 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1666464484
transform 1 0 5244 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1666464484
transform 1 0 8004 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1666464484
transform 1 0 10764 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1666464484
transform 1 0 13524 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1666464484
transform 1 0 16284 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1666464484
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1666464484
transform 1 0 21804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1666464484
transform 1 0 24564 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1666464484
transform 1 0 27324 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1666464484
transform 1 0 30084 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1666464484
transform 1 0 32844 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1666464484
transform 1 0 35604 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1666464484
transform 1 0 38364 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1666464484
transform 1 0 41124 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1666464484
transform 1 0 43884 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1666464484
transform 1 0 46644 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1666464484
transform 1 0 49404 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1666464484
transform 1 0 52164 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1666464484
transform 1 0 54924 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1666464484
transform 1 0 57684 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1666464484
transform 1 0 3864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1666464484
transform 1 0 6624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1666464484
transform 1 0 9384 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1666464484
transform 1 0 12144 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1666464484
transform 1 0 14904 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1666464484
transform 1 0 17664 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1666464484
transform 1 0 20424 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1666464484
transform 1 0 23184 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1666464484
transform 1 0 25944 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1666464484
transform 1 0 28704 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1666464484
transform 1 0 31464 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1666464484
transform 1 0 34224 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1666464484
transform 1 0 36984 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1666464484
transform 1 0 39744 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1666464484
transform 1 0 42504 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1666464484
transform 1 0 45264 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1666464484
transform 1 0 48024 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1666464484
transform 1 0 50784 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1666464484
transform 1 0 53544 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1666464484
transform 1 0 56304 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1666464484
transform 1 0 2484 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1666464484
transform 1 0 5244 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1666464484
transform 1 0 8004 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1666464484
transform 1 0 10764 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1666464484
transform 1 0 13524 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1666464484
transform 1 0 16284 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1666464484
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1666464484
transform 1 0 21804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1666464484
transform 1 0 24564 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1666464484
transform 1 0 27324 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1666464484
transform 1 0 30084 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1666464484
transform 1 0 32844 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1666464484
transform 1 0 35604 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1666464484
transform 1 0 38364 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1666464484
transform 1 0 41124 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1666464484
transform 1 0 43884 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1666464484
transform 1 0 46644 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1666464484
transform 1 0 49404 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1666464484
transform 1 0 52164 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1637
timestamp 1666464484
transform 1 0 54924 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1638
timestamp 1666464484
transform 1 0 57684 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1639
timestamp 1666464484
transform 1 0 3864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1640
timestamp 1666464484
transform 1 0 6624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1641
timestamp 1666464484
transform 1 0 9384 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1642
timestamp 1666464484
transform 1 0 12144 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1643
timestamp 1666464484
transform 1 0 14904 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1644
timestamp 1666464484
transform 1 0 17664 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1645
timestamp 1666464484
transform 1 0 20424 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1646
timestamp 1666464484
transform 1 0 23184 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1647
timestamp 1666464484
transform 1 0 25944 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1648
timestamp 1666464484
transform 1 0 28704 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1649
timestamp 1666464484
transform 1 0 31464 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1650
timestamp 1666464484
transform 1 0 34224 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1651
timestamp 1666464484
transform 1 0 36984 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1652
timestamp 1666464484
transform 1 0 39744 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1653
timestamp 1666464484
transform 1 0 42504 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1654
timestamp 1666464484
transform 1 0 45264 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1655
timestamp 1666464484
transform 1 0 48024 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1656
timestamp 1666464484
transform 1 0 50784 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1657
timestamp 1666464484
transform 1 0 53544 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1658
timestamp 1666464484
transform 1 0 56304 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1659
timestamp 1666464484
transform 1 0 2484 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1660
timestamp 1666464484
transform 1 0 5244 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1661
timestamp 1666464484
transform 1 0 8004 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1662
timestamp 1666464484
transform 1 0 10764 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1663
timestamp 1666464484
transform 1 0 13524 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1664
timestamp 1666464484
transform 1 0 16284 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1665
timestamp 1666464484
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1666
timestamp 1666464484
transform 1 0 21804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1667
timestamp 1666464484
transform 1 0 24564 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1668
timestamp 1666464484
transform 1 0 27324 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1669
timestamp 1666464484
transform 1 0 30084 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1670
timestamp 1666464484
transform 1 0 32844 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1671
timestamp 1666464484
transform 1 0 35604 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1672
timestamp 1666464484
transform 1 0 38364 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1673
timestamp 1666464484
transform 1 0 41124 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1674
timestamp 1666464484
transform 1 0 43884 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1675
timestamp 1666464484
transform 1 0 46644 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1676
timestamp 1666464484
transform 1 0 49404 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1677
timestamp 1666464484
transform 1 0 52164 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1678
timestamp 1666464484
transform 1 0 54924 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1679
timestamp 1666464484
transform 1 0 57684 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1680
timestamp 1666464484
transform 1 0 3864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1681
timestamp 1666464484
transform 1 0 6624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1682
timestamp 1666464484
transform 1 0 9384 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1683
timestamp 1666464484
transform 1 0 12144 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1684
timestamp 1666464484
transform 1 0 14904 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1685
timestamp 1666464484
transform 1 0 17664 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1686
timestamp 1666464484
transform 1 0 20424 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1687
timestamp 1666464484
transform 1 0 23184 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1688
timestamp 1666464484
transform 1 0 25944 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1689
timestamp 1666464484
transform 1 0 28704 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1690
timestamp 1666464484
transform 1 0 31464 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1691
timestamp 1666464484
transform 1 0 34224 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1692
timestamp 1666464484
transform 1 0 36984 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1693
timestamp 1666464484
transform 1 0 39744 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1694
timestamp 1666464484
transform 1 0 42504 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1695
timestamp 1666464484
transform 1 0 45264 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1696
timestamp 1666464484
transform 1 0 48024 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1697
timestamp 1666464484
transform 1 0 50784 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1698
timestamp 1666464484
transform 1 0 53544 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1699
timestamp 1666464484
transform 1 0 56304 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1700
timestamp 1666464484
transform 1 0 2484 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1701
timestamp 1666464484
transform 1 0 5244 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1702
timestamp 1666464484
transform 1 0 8004 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1703
timestamp 1666464484
transform 1 0 10764 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1704
timestamp 1666464484
transform 1 0 13524 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1705
timestamp 1666464484
transform 1 0 16284 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1706
timestamp 1666464484
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1707
timestamp 1666464484
transform 1 0 21804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1708
timestamp 1666464484
transform 1 0 24564 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1709
timestamp 1666464484
transform 1 0 27324 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1710
timestamp 1666464484
transform 1 0 30084 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1711
timestamp 1666464484
transform 1 0 32844 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1712
timestamp 1666464484
transform 1 0 35604 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1713
timestamp 1666464484
transform 1 0 38364 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1714
timestamp 1666464484
transform 1 0 41124 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1715
timestamp 1666464484
transform 1 0 43884 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1716
timestamp 1666464484
transform 1 0 46644 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1717
timestamp 1666464484
transform 1 0 49404 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1718
timestamp 1666464484
transform 1 0 52164 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1719
timestamp 1666464484
transform 1 0 54924 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1720
timestamp 1666464484
transform 1 0 57684 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1721
timestamp 1666464484
transform 1 0 3864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1722
timestamp 1666464484
transform 1 0 6624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1723
timestamp 1666464484
transform 1 0 9384 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1724
timestamp 1666464484
transform 1 0 12144 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1725
timestamp 1666464484
transform 1 0 14904 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1726
timestamp 1666464484
transform 1 0 17664 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1727
timestamp 1666464484
transform 1 0 20424 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1728
timestamp 1666464484
transform 1 0 23184 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1729
timestamp 1666464484
transform 1 0 25944 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1730
timestamp 1666464484
transform 1 0 28704 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1731
timestamp 1666464484
transform 1 0 31464 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1732
timestamp 1666464484
transform 1 0 34224 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1733
timestamp 1666464484
transform 1 0 36984 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1734
timestamp 1666464484
transform 1 0 39744 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1735
timestamp 1666464484
transform 1 0 42504 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1736
timestamp 1666464484
transform 1 0 45264 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1737
timestamp 1666464484
transform 1 0 48024 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1738
timestamp 1666464484
transform 1 0 50784 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1739
timestamp 1666464484
transform 1 0 53544 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1740
timestamp 1666464484
transform 1 0 56304 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1741
timestamp 1666464484
transform 1 0 2484 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1742
timestamp 1666464484
transform 1 0 5244 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1743
timestamp 1666464484
transform 1 0 8004 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1744
timestamp 1666464484
transform 1 0 10764 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1745
timestamp 1666464484
transform 1 0 13524 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1746
timestamp 1666464484
transform 1 0 16284 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1747
timestamp 1666464484
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1748
timestamp 1666464484
transform 1 0 21804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1749
timestamp 1666464484
transform 1 0 24564 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1750
timestamp 1666464484
transform 1 0 27324 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1751
timestamp 1666464484
transform 1 0 30084 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1752
timestamp 1666464484
transform 1 0 32844 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1753
timestamp 1666464484
transform 1 0 35604 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1754
timestamp 1666464484
transform 1 0 38364 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1755
timestamp 1666464484
transform 1 0 41124 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1756
timestamp 1666464484
transform 1 0 43884 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1757
timestamp 1666464484
transform 1 0 46644 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1758
timestamp 1666464484
transform 1 0 49404 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1759
timestamp 1666464484
transform 1 0 52164 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1760
timestamp 1666464484
transform 1 0 54924 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1761
timestamp 1666464484
transform 1 0 57684 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1762
timestamp 1666464484
transform 1 0 3864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1763
timestamp 1666464484
transform 1 0 6624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1764
timestamp 1666464484
transform 1 0 9384 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1765
timestamp 1666464484
transform 1 0 12144 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1766
timestamp 1666464484
transform 1 0 14904 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1767
timestamp 1666464484
transform 1 0 17664 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1768
timestamp 1666464484
transform 1 0 20424 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1769
timestamp 1666464484
transform 1 0 23184 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1770
timestamp 1666464484
transform 1 0 25944 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1771
timestamp 1666464484
transform 1 0 28704 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1772
timestamp 1666464484
transform 1 0 31464 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1773
timestamp 1666464484
transform 1 0 34224 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1774
timestamp 1666464484
transform 1 0 36984 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1775
timestamp 1666464484
transform 1 0 39744 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1776
timestamp 1666464484
transform 1 0 42504 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1777
timestamp 1666464484
transform 1 0 45264 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1778
timestamp 1666464484
transform 1 0 48024 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1779
timestamp 1666464484
transform 1 0 50784 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1780
timestamp 1666464484
transform 1 0 53544 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1781
timestamp 1666464484
transform 1 0 56304 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1782
timestamp 1666464484
transform 1 0 2484 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1783
timestamp 1666464484
transform 1 0 5244 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1784
timestamp 1666464484
transform 1 0 8004 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1785
timestamp 1666464484
transform 1 0 10764 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1786
timestamp 1666464484
transform 1 0 13524 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1787
timestamp 1666464484
transform 1 0 16284 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1788
timestamp 1666464484
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1789
timestamp 1666464484
transform 1 0 21804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1790
timestamp 1666464484
transform 1 0 24564 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1791
timestamp 1666464484
transform 1 0 27324 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1792
timestamp 1666464484
transform 1 0 30084 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1793
timestamp 1666464484
transform 1 0 32844 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1794
timestamp 1666464484
transform 1 0 35604 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1795
timestamp 1666464484
transform 1 0 38364 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1796
timestamp 1666464484
transform 1 0 41124 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1797
timestamp 1666464484
transform 1 0 43884 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1798
timestamp 1666464484
transform 1 0 46644 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1799
timestamp 1666464484
transform 1 0 49404 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1800
timestamp 1666464484
transform 1 0 52164 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1801
timestamp 1666464484
transform 1 0 54924 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1802
timestamp 1666464484
transform 1 0 57684 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1803
timestamp 1666464484
transform 1 0 3864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1804
timestamp 1666464484
transform 1 0 6624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1805
timestamp 1666464484
transform 1 0 9384 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1806
timestamp 1666464484
transform 1 0 12144 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1807
timestamp 1666464484
transform 1 0 14904 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1808
timestamp 1666464484
transform 1 0 17664 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1809
timestamp 1666464484
transform 1 0 20424 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1810
timestamp 1666464484
transform 1 0 23184 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1811
timestamp 1666464484
transform 1 0 25944 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1812
timestamp 1666464484
transform 1 0 28704 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1813
timestamp 1666464484
transform 1 0 31464 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1814
timestamp 1666464484
transform 1 0 34224 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1815
timestamp 1666464484
transform 1 0 36984 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1816
timestamp 1666464484
transform 1 0 39744 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1817
timestamp 1666464484
transform 1 0 42504 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1818
timestamp 1666464484
transform 1 0 45264 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1819
timestamp 1666464484
transform 1 0 48024 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1820
timestamp 1666464484
transform 1 0 50784 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1821
timestamp 1666464484
transform 1 0 53544 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1822
timestamp 1666464484
transform 1 0 56304 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1823
timestamp 1666464484
transform 1 0 2484 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1824
timestamp 1666464484
transform 1 0 5244 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1825
timestamp 1666464484
transform 1 0 8004 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1826
timestamp 1666464484
transform 1 0 10764 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1827
timestamp 1666464484
transform 1 0 13524 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1828
timestamp 1666464484
transform 1 0 16284 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1829
timestamp 1666464484
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1830
timestamp 1666464484
transform 1 0 21804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1831
timestamp 1666464484
transform 1 0 24564 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1832
timestamp 1666464484
transform 1 0 27324 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1833
timestamp 1666464484
transform 1 0 30084 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1834
timestamp 1666464484
transform 1 0 32844 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1835
timestamp 1666464484
transform 1 0 35604 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1836
timestamp 1666464484
transform 1 0 38364 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1837
timestamp 1666464484
transform 1 0 41124 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1838
timestamp 1666464484
transform 1 0 43884 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1839
timestamp 1666464484
transform 1 0 46644 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1840
timestamp 1666464484
transform 1 0 49404 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1841
timestamp 1666464484
transform 1 0 52164 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1842
timestamp 1666464484
transform 1 0 54924 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1843
timestamp 1666464484
transform 1 0 57684 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1844
timestamp 1666464484
transform 1 0 3864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1845
timestamp 1666464484
transform 1 0 6624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1846
timestamp 1666464484
transform 1 0 9384 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1847
timestamp 1666464484
transform 1 0 12144 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1848
timestamp 1666464484
transform 1 0 14904 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1849
timestamp 1666464484
transform 1 0 17664 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1850
timestamp 1666464484
transform 1 0 20424 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1851
timestamp 1666464484
transform 1 0 23184 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1852
timestamp 1666464484
transform 1 0 25944 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1853
timestamp 1666464484
transform 1 0 28704 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1854
timestamp 1666464484
transform 1 0 31464 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1855
timestamp 1666464484
transform 1 0 34224 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1856
timestamp 1666464484
transform 1 0 36984 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1857
timestamp 1666464484
transform 1 0 39744 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1858
timestamp 1666464484
transform 1 0 42504 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1859
timestamp 1666464484
transform 1 0 45264 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1860
timestamp 1666464484
transform 1 0 48024 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1861
timestamp 1666464484
transform 1 0 50784 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1862
timestamp 1666464484
transform 1 0 53544 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1863
timestamp 1666464484
transform 1 0 56304 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1864
timestamp 1666464484
transform 1 0 2484 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1865
timestamp 1666464484
transform 1 0 5244 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1866
timestamp 1666464484
transform 1 0 8004 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1867
timestamp 1666464484
transform 1 0 10764 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1868
timestamp 1666464484
transform 1 0 13524 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1869
timestamp 1666464484
transform 1 0 16284 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1870
timestamp 1666464484
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1871
timestamp 1666464484
transform 1 0 21804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1872
timestamp 1666464484
transform 1 0 24564 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1873
timestamp 1666464484
transform 1 0 27324 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1874
timestamp 1666464484
transform 1 0 30084 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1875
timestamp 1666464484
transform 1 0 32844 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1876
timestamp 1666464484
transform 1 0 35604 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1877
timestamp 1666464484
transform 1 0 38364 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1878
timestamp 1666464484
transform 1 0 41124 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1879
timestamp 1666464484
transform 1 0 43884 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1880
timestamp 1666464484
transform 1 0 46644 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1881
timestamp 1666464484
transform 1 0 49404 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1882
timestamp 1666464484
transform 1 0 52164 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1883
timestamp 1666464484
transform 1 0 54924 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1884
timestamp 1666464484
transform 1 0 57684 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1885
timestamp 1666464484
transform 1 0 3864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1886
timestamp 1666464484
transform 1 0 6624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1887
timestamp 1666464484
transform 1 0 9384 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1888
timestamp 1666464484
transform 1 0 12144 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1889
timestamp 1666464484
transform 1 0 14904 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1890
timestamp 1666464484
transform 1 0 17664 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1891
timestamp 1666464484
transform 1 0 20424 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1892
timestamp 1666464484
transform 1 0 23184 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1893
timestamp 1666464484
transform 1 0 25944 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1894
timestamp 1666464484
transform 1 0 28704 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1895
timestamp 1666464484
transform 1 0 31464 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1896
timestamp 1666464484
transform 1 0 34224 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1897
timestamp 1666464484
transform 1 0 36984 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1898
timestamp 1666464484
transform 1 0 39744 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1899
timestamp 1666464484
transform 1 0 42504 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1900
timestamp 1666464484
transform 1 0 45264 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1901
timestamp 1666464484
transform 1 0 48024 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1902
timestamp 1666464484
transform 1 0 50784 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1903
timestamp 1666464484
transform 1 0 53544 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1904
timestamp 1666464484
transform 1 0 56304 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1905
timestamp 1666464484
transform 1 0 2484 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1906
timestamp 1666464484
transform 1 0 5244 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1907
timestamp 1666464484
transform 1 0 8004 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1908
timestamp 1666464484
transform 1 0 10764 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1909
timestamp 1666464484
transform 1 0 13524 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1910
timestamp 1666464484
transform 1 0 16284 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1911
timestamp 1666464484
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1912
timestamp 1666464484
transform 1 0 21804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1913
timestamp 1666464484
transform 1 0 24564 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1914
timestamp 1666464484
transform 1 0 27324 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1915
timestamp 1666464484
transform 1 0 30084 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1916
timestamp 1666464484
transform 1 0 32844 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1917
timestamp 1666464484
transform 1 0 35604 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1918
timestamp 1666464484
transform 1 0 38364 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1919
timestamp 1666464484
transform 1 0 41124 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1920
timestamp 1666464484
transform 1 0 43884 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1921
timestamp 1666464484
transform 1 0 46644 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1922
timestamp 1666464484
transform 1 0 49404 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1923
timestamp 1666464484
transform 1 0 52164 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1924
timestamp 1666464484
transform 1 0 54924 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1925
timestamp 1666464484
transform 1 0 57684 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1926
timestamp 1666464484
transform 1 0 3864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1927
timestamp 1666464484
transform 1 0 6624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1928
timestamp 1666464484
transform 1 0 9384 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1929
timestamp 1666464484
transform 1 0 12144 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1930
timestamp 1666464484
transform 1 0 14904 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1931
timestamp 1666464484
transform 1 0 17664 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1932
timestamp 1666464484
transform 1 0 20424 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1933
timestamp 1666464484
transform 1 0 23184 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1934
timestamp 1666464484
transform 1 0 25944 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1935
timestamp 1666464484
transform 1 0 28704 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1936
timestamp 1666464484
transform 1 0 31464 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1937
timestamp 1666464484
transform 1 0 34224 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1938
timestamp 1666464484
transform 1 0 36984 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1939
timestamp 1666464484
transform 1 0 39744 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1940
timestamp 1666464484
transform 1 0 42504 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1941
timestamp 1666464484
transform 1 0 45264 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1942
timestamp 1666464484
transform 1 0 48024 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1943
timestamp 1666464484
transform 1 0 50784 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1944
timestamp 1666464484
transform 1 0 53544 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1945
timestamp 1666464484
transform 1 0 56304 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1946
timestamp 1666464484
transform 1 0 2484 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1947
timestamp 1666464484
transform 1 0 5244 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1948
timestamp 1666464484
transform 1 0 8004 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1949
timestamp 1666464484
transform 1 0 10764 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1950
timestamp 1666464484
transform 1 0 13524 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1951
timestamp 1666464484
transform 1 0 16284 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1952
timestamp 1666464484
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1953
timestamp 1666464484
transform 1 0 21804 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1954
timestamp 1666464484
transform 1 0 24564 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1955
timestamp 1666464484
transform 1 0 27324 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1956
timestamp 1666464484
transform 1 0 30084 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1957
timestamp 1666464484
transform 1 0 32844 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1958
timestamp 1666464484
transform 1 0 35604 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1959
timestamp 1666464484
transform 1 0 38364 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1960
timestamp 1666464484
transform 1 0 41124 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1961
timestamp 1666464484
transform 1 0 43884 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1962
timestamp 1666464484
transform 1 0 46644 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1963
timestamp 1666464484
transform 1 0 49404 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1964
timestamp 1666464484
transform 1 0 52164 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1965
timestamp 1666464484
transform 1 0 54924 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1966
timestamp 1666464484
transform 1 0 57684 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1967
timestamp 1666464484
transform 1 0 3864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1968
timestamp 1666464484
transform 1 0 6624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1969
timestamp 1666464484
transform 1 0 9384 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1970
timestamp 1666464484
transform 1 0 12144 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1971
timestamp 1666464484
transform 1 0 14904 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1972
timestamp 1666464484
transform 1 0 17664 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1973
timestamp 1666464484
transform 1 0 20424 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1974
timestamp 1666464484
transform 1 0 23184 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1975
timestamp 1666464484
transform 1 0 25944 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1976
timestamp 1666464484
transform 1 0 28704 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1977
timestamp 1666464484
transform 1 0 31464 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1978
timestamp 1666464484
transform 1 0 34224 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1979
timestamp 1666464484
transform 1 0 36984 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1980
timestamp 1666464484
transform 1 0 39744 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1981
timestamp 1666464484
transform 1 0 42504 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1982
timestamp 1666464484
transform 1 0 45264 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1983
timestamp 1666464484
transform 1 0 48024 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1984
timestamp 1666464484
transform 1 0 50784 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1985
timestamp 1666464484
transform 1 0 53544 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1986
timestamp 1666464484
transform 1 0 56304 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1987
timestamp 1666464484
transform 1 0 2484 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1988
timestamp 1666464484
transform 1 0 5244 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1989
timestamp 1666464484
transform 1 0 8004 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1990
timestamp 1666464484
transform 1 0 10764 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1991
timestamp 1666464484
transform 1 0 13524 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1992
timestamp 1666464484
transform 1 0 16284 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1993
timestamp 1666464484
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1994
timestamp 1666464484
transform 1 0 21804 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1995
timestamp 1666464484
transform 1 0 24564 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1996
timestamp 1666464484
transform 1 0 27324 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1997
timestamp 1666464484
transform 1 0 30084 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1998
timestamp 1666464484
transform 1 0 32844 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1999
timestamp 1666464484
transform 1 0 35604 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2000
timestamp 1666464484
transform 1 0 38364 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2001
timestamp 1666464484
transform 1 0 41124 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2002
timestamp 1666464484
transform 1 0 43884 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2003
timestamp 1666464484
transform 1 0 46644 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2004
timestamp 1666464484
transform 1 0 49404 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2005
timestamp 1666464484
transform 1 0 52164 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2006
timestamp 1666464484
transform 1 0 54924 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2007
timestamp 1666464484
transform 1 0 57684 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2008
timestamp 1666464484
transform 1 0 3864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2009
timestamp 1666464484
transform 1 0 6624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2010
timestamp 1666464484
transform 1 0 9384 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2011
timestamp 1666464484
transform 1 0 12144 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2012
timestamp 1666464484
transform 1 0 14904 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2013
timestamp 1666464484
transform 1 0 17664 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2014
timestamp 1666464484
transform 1 0 20424 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2015
timestamp 1666464484
transform 1 0 23184 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2016
timestamp 1666464484
transform 1 0 25944 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2017
timestamp 1666464484
transform 1 0 28704 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2018
timestamp 1666464484
transform 1 0 31464 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2019
timestamp 1666464484
transform 1 0 34224 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2020
timestamp 1666464484
transform 1 0 36984 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2021
timestamp 1666464484
transform 1 0 39744 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2022
timestamp 1666464484
transform 1 0 42504 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2023
timestamp 1666464484
transform 1 0 45264 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2024
timestamp 1666464484
transform 1 0 48024 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2025
timestamp 1666464484
transform 1 0 50784 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2026
timestamp 1666464484
transform 1 0 53544 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2027
timestamp 1666464484
transform 1 0 56304 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2028
timestamp 1666464484
transform 1 0 2484 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2029
timestamp 1666464484
transform 1 0 5244 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2030
timestamp 1666464484
transform 1 0 8004 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2031
timestamp 1666464484
transform 1 0 10764 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2032
timestamp 1666464484
transform 1 0 13524 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2033
timestamp 1666464484
transform 1 0 16284 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2034
timestamp 1666464484
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2035
timestamp 1666464484
transform 1 0 21804 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2036
timestamp 1666464484
transform 1 0 24564 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2037
timestamp 1666464484
transform 1 0 27324 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2038
timestamp 1666464484
transform 1 0 30084 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2039
timestamp 1666464484
transform 1 0 32844 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2040
timestamp 1666464484
transform 1 0 35604 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2041
timestamp 1666464484
transform 1 0 38364 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2042
timestamp 1666464484
transform 1 0 41124 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2043
timestamp 1666464484
transform 1 0 43884 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2044
timestamp 1666464484
transform 1 0 46644 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2045
timestamp 1666464484
transform 1 0 49404 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2046
timestamp 1666464484
transform 1 0 52164 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2047
timestamp 1666464484
transform 1 0 54924 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2048
timestamp 1666464484
transform 1 0 57684 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2049
timestamp 1666464484
transform 1 0 3864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2050
timestamp 1666464484
transform 1 0 6624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2051
timestamp 1666464484
transform 1 0 9384 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2052
timestamp 1666464484
transform 1 0 12144 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2053
timestamp 1666464484
transform 1 0 14904 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2054
timestamp 1666464484
transform 1 0 17664 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2055
timestamp 1666464484
transform 1 0 20424 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2056
timestamp 1666464484
transform 1 0 23184 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2057
timestamp 1666464484
transform 1 0 25944 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2058
timestamp 1666464484
transform 1 0 28704 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2059
timestamp 1666464484
transform 1 0 31464 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2060
timestamp 1666464484
transform 1 0 34224 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2061
timestamp 1666464484
transform 1 0 36984 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2062
timestamp 1666464484
transform 1 0 39744 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2063
timestamp 1666464484
transform 1 0 42504 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2064
timestamp 1666464484
transform 1 0 45264 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2065
timestamp 1666464484
transform 1 0 48024 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2066
timestamp 1666464484
transform 1 0 50784 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2067
timestamp 1666464484
transform 1 0 53544 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2068
timestamp 1666464484
transform 1 0 56304 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2069
timestamp 1666464484
transform 1 0 2484 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2070
timestamp 1666464484
transform 1 0 5244 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2071
timestamp 1666464484
transform 1 0 8004 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2072
timestamp 1666464484
transform 1 0 10764 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2073
timestamp 1666464484
transform 1 0 13524 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2074
timestamp 1666464484
transform 1 0 16284 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2075
timestamp 1666464484
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2076
timestamp 1666464484
transform 1 0 21804 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2077
timestamp 1666464484
transform 1 0 24564 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2078
timestamp 1666464484
transform 1 0 27324 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2079
timestamp 1666464484
transform 1 0 30084 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2080
timestamp 1666464484
transform 1 0 32844 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2081
timestamp 1666464484
transform 1 0 35604 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2082
timestamp 1666464484
transform 1 0 38364 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2083
timestamp 1666464484
transform 1 0 41124 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2084
timestamp 1666464484
transform 1 0 43884 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2085
timestamp 1666464484
transform 1 0 46644 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2086
timestamp 1666464484
transform 1 0 49404 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2087
timestamp 1666464484
transform 1 0 52164 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2088
timestamp 1666464484
transform 1 0 54924 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2089
timestamp 1666464484
transform 1 0 57684 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2090
timestamp 1666464484
transform 1 0 3864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2091
timestamp 1666464484
transform 1 0 6624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2092
timestamp 1666464484
transform 1 0 9384 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2093
timestamp 1666464484
transform 1 0 12144 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2094
timestamp 1666464484
transform 1 0 14904 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2095
timestamp 1666464484
transform 1 0 17664 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2096
timestamp 1666464484
transform 1 0 20424 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2097
timestamp 1666464484
transform 1 0 23184 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2098
timestamp 1666464484
transform 1 0 25944 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2099
timestamp 1666464484
transform 1 0 28704 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2100
timestamp 1666464484
transform 1 0 31464 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2101
timestamp 1666464484
transform 1 0 34224 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2102
timestamp 1666464484
transform 1 0 36984 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2103
timestamp 1666464484
transform 1 0 39744 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2104
timestamp 1666464484
transform 1 0 42504 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2105
timestamp 1666464484
transform 1 0 45264 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2106
timestamp 1666464484
transform 1 0 48024 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2107
timestamp 1666464484
transform 1 0 50784 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2108
timestamp 1666464484
transform 1 0 53544 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2109
timestamp 1666464484
transform 1 0 56304 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2110
timestamp 1666464484
transform 1 0 2484 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2111
timestamp 1666464484
transform 1 0 5244 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2112
timestamp 1666464484
transform 1 0 8004 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2113
timestamp 1666464484
transform 1 0 10764 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2114
timestamp 1666464484
transform 1 0 13524 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2115
timestamp 1666464484
transform 1 0 16284 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2116
timestamp 1666464484
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2117
timestamp 1666464484
transform 1 0 21804 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2118
timestamp 1666464484
transform 1 0 24564 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2119
timestamp 1666464484
transform 1 0 27324 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2120
timestamp 1666464484
transform 1 0 30084 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2121
timestamp 1666464484
transform 1 0 32844 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2122
timestamp 1666464484
transform 1 0 35604 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2123
timestamp 1666464484
transform 1 0 38364 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2124
timestamp 1666464484
transform 1 0 41124 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2125
timestamp 1666464484
transform 1 0 43884 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2126
timestamp 1666464484
transform 1 0 46644 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2127
timestamp 1666464484
transform 1 0 49404 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2128
timestamp 1666464484
transform 1 0 52164 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2129
timestamp 1666464484
transform 1 0 54924 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2130
timestamp 1666464484
transform 1 0 57684 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2131
timestamp 1666464484
transform 1 0 3864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2132
timestamp 1666464484
transform 1 0 6624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2133
timestamp 1666464484
transform 1 0 9384 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2134
timestamp 1666464484
transform 1 0 12144 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2135
timestamp 1666464484
transform 1 0 14904 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2136
timestamp 1666464484
transform 1 0 17664 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2137
timestamp 1666464484
transform 1 0 20424 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2138
timestamp 1666464484
transform 1 0 23184 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2139
timestamp 1666464484
transform 1 0 25944 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2140
timestamp 1666464484
transform 1 0 28704 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2141
timestamp 1666464484
transform 1 0 31464 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2142
timestamp 1666464484
transform 1 0 34224 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2143
timestamp 1666464484
transform 1 0 36984 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2144
timestamp 1666464484
transform 1 0 39744 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2145
timestamp 1666464484
transform 1 0 42504 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2146
timestamp 1666464484
transform 1 0 45264 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2147
timestamp 1666464484
transform 1 0 48024 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2148
timestamp 1666464484
transform 1 0 50784 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2149
timestamp 1666464484
transform 1 0 53544 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2150
timestamp 1666464484
transform 1 0 56304 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2151
timestamp 1666464484
transform 1 0 2484 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2152
timestamp 1666464484
transform 1 0 5244 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2153
timestamp 1666464484
transform 1 0 8004 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2154
timestamp 1666464484
transform 1 0 10764 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2155
timestamp 1666464484
transform 1 0 13524 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2156
timestamp 1666464484
transform 1 0 16284 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2157
timestamp 1666464484
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2158
timestamp 1666464484
transform 1 0 21804 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2159
timestamp 1666464484
transform 1 0 24564 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2160
timestamp 1666464484
transform 1 0 27324 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2161
timestamp 1666464484
transform 1 0 30084 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2162
timestamp 1666464484
transform 1 0 32844 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2163
timestamp 1666464484
transform 1 0 35604 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2164
timestamp 1666464484
transform 1 0 38364 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2165
timestamp 1666464484
transform 1 0 41124 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2166
timestamp 1666464484
transform 1 0 43884 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2167
timestamp 1666464484
transform 1 0 46644 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2168
timestamp 1666464484
transform 1 0 49404 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2169
timestamp 1666464484
transform 1 0 52164 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2170
timestamp 1666464484
transform 1 0 54924 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2171
timestamp 1666464484
transform 1 0 57684 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2172
timestamp 1666464484
transform 1 0 3864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2173
timestamp 1666464484
transform 1 0 6624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2174
timestamp 1666464484
transform 1 0 9384 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2175
timestamp 1666464484
transform 1 0 12144 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2176
timestamp 1666464484
transform 1 0 14904 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2177
timestamp 1666464484
transform 1 0 17664 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2178
timestamp 1666464484
transform 1 0 20424 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2179
timestamp 1666464484
transform 1 0 23184 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2180
timestamp 1666464484
transform 1 0 25944 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2181
timestamp 1666464484
transform 1 0 28704 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2182
timestamp 1666464484
transform 1 0 31464 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2183
timestamp 1666464484
transform 1 0 34224 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2184
timestamp 1666464484
transform 1 0 36984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2185
timestamp 1666464484
transform 1 0 39744 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2186
timestamp 1666464484
transform 1 0 42504 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2187
timestamp 1666464484
transform 1 0 45264 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2188
timestamp 1666464484
transform 1 0 48024 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2189
timestamp 1666464484
transform 1 0 50784 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2190
timestamp 1666464484
transform 1 0 53544 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2191
timestamp 1666464484
transform 1 0 56304 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2192
timestamp 1666464484
transform 1 0 2484 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2193
timestamp 1666464484
transform 1 0 5244 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2194
timestamp 1666464484
transform 1 0 8004 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2195
timestamp 1666464484
transform 1 0 10764 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2196
timestamp 1666464484
transform 1 0 13524 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2197
timestamp 1666464484
transform 1 0 16284 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2198
timestamp 1666464484
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2199
timestamp 1666464484
transform 1 0 21804 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2200
timestamp 1666464484
transform 1 0 24564 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2201
timestamp 1666464484
transform 1 0 27324 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2202
timestamp 1666464484
transform 1 0 30084 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2203
timestamp 1666464484
transform 1 0 32844 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2204
timestamp 1666464484
transform 1 0 35604 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2205
timestamp 1666464484
transform 1 0 38364 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2206
timestamp 1666464484
transform 1 0 41124 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2207
timestamp 1666464484
transform 1 0 43884 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2208
timestamp 1666464484
transform 1 0 46644 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2209
timestamp 1666464484
transform 1 0 49404 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2210
timestamp 1666464484
transform 1 0 52164 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2211
timestamp 1666464484
transform 1 0 54924 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2212
timestamp 1666464484
transform 1 0 57684 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2213
timestamp 1666464484
transform 1 0 3864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2214
timestamp 1666464484
transform 1 0 6624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2215
timestamp 1666464484
transform 1 0 9384 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2216
timestamp 1666464484
transform 1 0 12144 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2217
timestamp 1666464484
transform 1 0 14904 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2218
timestamp 1666464484
transform 1 0 17664 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2219
timestamp 1666464484
transform 1 0 20424 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2220
timestamp 1666464484
transform 1 0 23184 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2221
timestamp 1666464484
transform 1 0 25944 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2222
timestamp 1666464484
transform 1 0 28704 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2223
timestamp 1666464484
transform 1 0 31464 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2224
timestamp 1666464484
transform 1 0 34224 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2225
timestamp 1666464484
transform 1 0 36984 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2226
timestamp 1666464484
transform 1 0 39744 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2227
timestamp 1666464484
transform 1 0 42504 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2228
timestamp 1666464484
transform 1 0 45264 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2229
timestamp 1666464484
transform 1 0 48024 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2230
timestamp 1666464484
transform 1 0 50784 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2231
timestamp 1666464484
transform 1 0 53544 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2232
timestamp 1666464484
transform 1 0 56304 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2233
timestamp 1666464484
transform 1 0 2484 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2234
timestamp 1666464484
transform 1 0 5244 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2235
timestamp 1666464484
transform 1 0 8004 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2236
timestamp 1666464484
transform 1 0 10764 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2237
timestamp 1666464484
transform 1 0 13524 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2238
timestamp 1666464484
transform 1 0 16284 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2239
timestamp 1666464484
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2240
timestamp 1666464484
transform 1 0 21804 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2241
timestamp 1666464484
transform 1 0 24564 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2242
timestamp 1666464484
transform 1 0 27324 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2243
timestamp 1666464484
transform 1 0 30084 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2244
timestamp 1666464484
transform 1 0 32844 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2245
timestamp 1666464484
transform 1 0 35604 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2246
timestamp 1666464484
transform 1 0 38364 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2247
timestamp 1666464484
transform 1 0 41124 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2248
timestamp 1666464484
transform 1 0 43884 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2249
timestamp 1666464484
transform 1 0 46644 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2250
timestamp 1666464484
transform 1 0 49404 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2251
timestamp 1666464484
transform 1 0 52164 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2252
timestamp 1666464484
transform 1 0 54924 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2253
timestamp 1666464484
transform 1 0 57684 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2254
timestamp 1666464484
transform 1 0 3864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2255
timestamp 1666464484
transform 1 0 6624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2256
timestamp 1666464484
transform 1 0 9384 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2257
timestamp 1666464484
transform 1 0 12144 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2258
timestamp 1666464484
transform 1 0 14904 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2259
timestamp 1666464484
transform 1 0 17664 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2260
timestamp 1666464484
transform 1 0 20424 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2261
timestamp 1666464484
transform 1 0 23184 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2262
timestamp 1666464484
transform 1 0 25944 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2263
timestamp 1666464484
transform 1 0 28704 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2264
timestamp 1666464484
transform 1 0 31464 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2265
timestamp 1666464484
transform 1 0 34224 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2266
timestamp 1666464484
transform 1 0 36984 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2267
timestamp 1666464484
transform 1 0 39744 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2268
timestamp 1666464484
transform 1 0 42504 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2269
timestamp 1666464484
transform 1 0 45264 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2270
timestamp 1666464484
transform 1 0 48024 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2271
timestamp 1666464484
transform 1 0 50784 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2272
timestamp 1666464484
transform 1 0 53544 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2273
timestamp 1666464484
transform 1 0 56304 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2274
timestamp 1666464484
transform 1 0 2484 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2275
timestamp 1666464484
transform 1 0 5244 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2276
timestamp 1666464484
transform 1 0 8004 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2277
timestamp 1666464484
transform 1 0 10764 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2278
timestamp 1666464484
transform 1 0 13524 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2279
timestamp 1666464484
transform 1 0 16284 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2280
timestamp 1666464484
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2281
timestamp 1666464484
transform 1 0 21804 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2282
timestamp 1666464484
transform 1 0 24564 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2283
timestamp 1666464484
transform 1 0 27324 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2284
timestamp 1666464484
transform 1 0 30084 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2285
timestamp 1666464484
transform 1 0 32844 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2286
timestamp 1666464484
transform 1 0 35604 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2287
timestamp 1666464484
transform 1 0 38364 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2288
timestamp 1666464484
transform 1 0 41124 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2289
timestamp 1666464484
transform 1 0 43884 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2290
timestamp 1666464484
transform 1 0 46644 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2291
timestamp 1666464484
transform 1 0 49404 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2292
timestamp 1666464484
transform 1 0 52164 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2293
timestamp 1666464484
transform 1 0 54924 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2294
timestamp 1666464484
transform 1 0 57684 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2295
timestamp 1666464484
transform 1 0 2484 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2296
timestamp 1666464484
transform 1 0 3864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2297
timestamp 1666464484
transform 1 0 5244 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2298
timestamp 1666464484
transform 1 0 6624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2299
timestamp 1666464484
transform 1 0 8004 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2300
timestamp 1666464484
transform 1 0 9384 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2301
timestamp 1666464484
transform 1 0 10764 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2302
timestamp 1666464484
transform 1 0 12144 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2303
timestamp 1666464484
transform 1 0 13524 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2304
timestamp 1666464484
transform 1 0 14904 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2305
timestamp 1666464484
transform 1 0 16284 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2306
timestamp 1666464484
transform 1 0 17664 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2307
timestamp 1666464484
transform 1 0 19044 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2308
timestamp 1666464484
transform 1 0 20424 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2309
timestamp 1666464484
transform 1 0 21804 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2310
timestamp 1666464484
transform 1 0 23184 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2311
timestamp 1666464484
transform 1 0 24564 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2312
timestamp 1666464484
transform 1 0 25944 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2313
timestamp 1666464484
transform 1 0 27324 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2314
timestamp 1666464484
transform 1 0 28704 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2315
timestamp 1666464484
transform 1 0 30084 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2316
timestamp 1666464484
transform 1 0 31464 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2317
timestamp 1666464484
transform 1 0 32844 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2318
timestamp 1666464484
transform 1 0 34224 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2319
timestamp 1666464484
transform 1 0 35604 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2320
timestamp 1666464484
transform 1 0 36984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2321
timestamp 1666464484
transform 1 0 38364 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2322
timestamp 1666464484
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2323
timestamp 1666464484
transform 1 0 41124 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2324
timestamp 1666464484
transform 1 0 42504 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2325
timestamp 1666464484
transform 1 0 43884 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2326
timestamp 1666464484
transform 1 0 45264 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2327
timestamp 1666464484
transform 1 0 46644 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2328
timestamp 1666464484
transform 1 0 48024 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2329
timestamp 1666464484
transform 1 0 49404 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2330
timestamp 1666464484
transform 1 0 50784 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2331
timestamp 1666464484
transform 1 0 52164 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2332
timestamp 1666464484
transform 1 0 53544 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2333
timestamp 1666464484
transform 1 0 54924 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2334
timestamp 1666464484
transform 1 0 56304 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2335
timestamp 1666464484
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _157_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27048 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _158_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _159_
timestamp 1666464484
transform 1 0 30820 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _160_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 37904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1666464484
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1666464484
transform -1 0 36800 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1666464484
transform 1 0 35880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1666464484
transform 1 0 34500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1666464484
transform 1 0 32660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1666464484
transform -1 0 35420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1666464484
transform -1 0 34040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1666464484
transform -1 0 33396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _170_
timestamp 1666464484
transform 1 0 31740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1666464484
transform 1 0 30728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1666464484
transform 1 0 32384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1666464484
transform 1 0 27600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1666464484
transform 1 0 29624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1666464484
transform 1 0 28244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1666464484
transform -1 0 30360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1666464484
transform -1 0 29716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1666464484
transform -1 0 29624 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1666464484
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1666464484
transform -1 0 25116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _181_
timestamp 1666464484
transform -1 0 25760 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1666464484
transform 1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1666464484
transform 1 0 22724 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1666464484
transform 1 0 24104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1666464484
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1666464484
transform 1 0 27324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1666464484
transform 1 0 26220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1666464484
transform -1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1666464484
transform 1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1666464484
transform -1 0 21712 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1666464484
transform -1 0 23092 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1666464484
transform -1 0 25760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _193_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 36340 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _194_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34500 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _195_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34776 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _196_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 28244 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _197_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 36432 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _198_
timestamp 1666464484
transform -1 0 35328 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _199_
timestamp 1666464484
transform -1 0 29624 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _200_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 35052 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _201_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34316 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _202_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32844 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _203_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31832 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _204_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 33580 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _205_
timestamp 1666464484
transform 1 0 31924 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _206_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30544 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _207_
timestamp 1666464484
transform -1 0 30452 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _208_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29072 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _209_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34500 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _210_
timestamp 1666464484
transform -1 0 27140 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _211_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28612 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _212_
timestamp 1666464484
transform -1 0 28520 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _213_
timestamp 1666464484
transform -1 0 44620 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _214_
timestamp 1666464484
transform 1 0 43792 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _215_
timestamp 1666464484
transform -1 0 43424 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _216_
timestamp 1666464484
transform 1 0 37720 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _217_
timestamp 1666464484
transform 1 0 43792 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _218_
timestamp 1666464484
transform -1 0 43424 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _219_
timestamp 1666464484
transform -1 0 39100 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _220_
timestamp 1666464484
transform -1 0 42872 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _221_
timestamp 1666464484
transform 1 0 41584 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _222_
timestamp 1666464484
transform 1 0 41400 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _223_
timestamp 1666464484
transform 1 0 40204 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _224_
timestamp 1666464484
transform -1 0 42228 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _225_
timestamp 1666464484
transform 1 0 40296 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _226_
timestamp 1666464484
transform 1 0 36800 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _227_
timestamp 1666464484
transform -1 0 38456 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _228_
timestamp 1666464484
transform -1 0 39284 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _229_
timestamp 1666464484
transform -1 0 43056 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _230_
timestamp 1666464484
transform -1 0 39560 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _231_
timestamp 1666464484
transform 1 0 38640 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _232_
timestamp 1666464484
transform -1 0 36800 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _233_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35236 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _234_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27968 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _235_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27600 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1666464484
transform -1 0 35420 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _237_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31740 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _238_
timestamp 1666464484
transform 1 0 31740 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _239_
timestamp 1666464484
transform 1 0 30728 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1666464484
transform -1 0 42320 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _241_
timestamp 1666464484
transform 1 0 40204 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _242_
timestamp 1666464484
transform -1 0 40572 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _243_
timestamp 1666464484
transform 1 0 40020 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _244_
timestamp 1666464484
transform -1 0 24472 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _245_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22264 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _246_
timestamp 1666464484
transform 1 0 23920 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1666464484
transform 1 0 24104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _248_
timestamp 1666464484
transform -1 0 24380 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _249_
timestamp 1666464484
transform -1 0 33304 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _250_
timestamp 1666464484
transform 1 0 32016 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _251_
timestamp 1666464484
transform 1 0 34500 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _252_
timestamp 1666464484
transform 1 0 33212 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _253_
timestamp 1666464484
transform 1 0 32660 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _254_
timestamp 1666464484
transform 1 0 40848 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _255_
timestamp 1666464484
transform -1 0 42044 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _256_
timestamp 1666464484
transform 1 0 42504 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _257_
timestamp 1666464484
transform 1 0 41492 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _258_
timestamp 1666464484
transform 1 0 41124 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _259_
timestamp 1666464484
transform 1 0 25300 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1666464484
transform 1 0 25484 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _261_
timestamp 1666464484
transform 1 0 25300 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1666464484
transform -1 0 25852 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _263_
timestamp 1666464484
transform 1 0 25116 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _264_
timestamp 1666464484
transform 1 0 31924 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _265_
timestamp 1666464484
transform 1 0 33120 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _266_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31004 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _267_
timestamp 1666464484
transform -1 0 31280 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _268_
timestamp 1666464484
transform -1 0 30452 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _269_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31556 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _270_
timestamp 1666464484
transform 1 0 41768 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _271_
timestamp 1666464484
transform 1 0 43240 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _272_
timestamp 1666464484
transform 1 0 38824 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _273_
timestamp 1666464484
transform 1 0 39468 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _274_
timestamp 1666464484
transform 1 0 40020 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _275_
timestamp 1666464484
transform -1 0 40756 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _276_
timestamp 1666464484
transform 1 0 26680 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1666464484
transform 1 0 26864 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _278_
timestamp 1666464484
transform -1 0 27600 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _279_
timestamp 1666464484
transform -1 0 25484 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _280_
timestamp 1666464484
transform -1 0 27140 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _281_
timestamp 1666464484
transform -1 0 29716 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _282_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27968 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _283_
timestamp 1666464484
transform 1 0 28612 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _284_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30820 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _285_
timestamp 1666464484
transform 1 0 33120 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _286_
timestamp 1666464484
transform 1 0 34224 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _287_
timestamp 1666464484
transform -1 0 28244 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _288_
timestamp 1666464484
transform 1 0 37628 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _289_
timestamp 1666464484
transform -1 0 38824 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _290_
timestamp 1666464484
transform -1 0 37904 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _291_
timestamp 1666464484
transform 1 0 44160 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _292_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 44160 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _293_
timestamp 1666464484
transform 1 0 37260 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _294_
timestamp 1666464484
transform 1 0 35972 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _295_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29900 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _296_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28980 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _519__194 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25208 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _520__195
timestamp 1666464484
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _520_
timestamp 1666464484
transform 1 0 22448 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _521_
timestamp 1666464484
transform 1 0 25208 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _521__196
timestamp 1666464484
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _522_
timestamp 1666464484
transform 1 0 23828 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _522__197
timestamp 1666464484
transform 1 0 22724 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _523__198
timestamp 1666464484
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _523_
timestamp 1666464484
transform 1 0 23828 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _524_
timestamp 1666464484
transform 1 0 26588 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _524__199
timestamp 1666464484
transform 1 0 23920 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _525__200
timestamp 1666464484
transform -1 0 27140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _525_
timestamp 1666464484
transform 1 0 26588 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _526__201
timestamp 1666464484
transform -1 0 27876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _526_
timestamp 1666464484
transform 1 0 27600 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _527__202
timestamp 1666464484
transform -1 0 28244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _527_
timestamp 1666464484
transform 1 0 27968 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _528_
timestamp 1666464484
transform 1 0 27876 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _528__203
timestamp 1666464484
transform 1 0 22724 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _529__204
timestamp 1666464484
transform 1 0 23460 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _529_
timestamp 1666464484
transform 1 0 25208 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _530_
timestamp 1666464484
transform 1 0 26588 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _530__205
timestamp 1666464484
transform 1 0 24104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _531_
timestamp 1666464484
transform 1 0 26588 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _531__206
timestamp 1666464484
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _532__207
timestamp 1666464484
transform 1 0 28244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _532_
timestamp 1666464484
transform 1 0 29164 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _533__208
timestamp 1666464484
transform 1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _533_
timestamp 1666464484
transform 1 0 29256 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _534__209
timestamp 1666464484
transform -1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _534_
timestamp 1666464484
transform 1 0 29348 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _535_
timestamp 1666464484
transform 1 0 30360 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _535__210
timestamp 1666464484
transform 1 0 28980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _536_
timestamp 1666464484
transform 1 0 30544 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _536__211
timestamp 1666464484
transform -1 0 30912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _537_
timestamp 1666464484
transform 1 0 29348 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _537__212
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _538__213
timestamp 1666464484
transform 1 0 32660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _538_
timestamp 1666464484
transform -1 0 33672 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _539__214
timestamp 1666464484
transform -1 0 32016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _539_
timestamp 1666464484
transform 1 0 30728 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _540_
timestamp 1666464484
transform -1 0 33672 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _540__215
timestamp 1666464484
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _541_
timestamp 1666464484
transform 1 0 33120 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _541__216
timestamp 1666464484
transform 1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _542_
timestamp 1666464484
transform 1 0 34500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _542__217
timestamp 1666464484
transform -1 0 34776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _543__218
timestamp 1666464484
transform -1 0 33580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _543_
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _544__219
timestamp 1666464484
transform -1 0 33396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _544_
timestamp 1666464484
transform 1 0 33120 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _545__220
timestamp 1666464484
transform 1 0 33764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _545_
timestamp 1666464484
transform -1 0 35052 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _546_
timestamp 1666464484
transform 1 0 35880 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _546__221
timestamp 1666464484
transform -1 0 36800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _547__222
timestamp 1666464484
transform 1 0 35880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _547_
timestamp 1666464484
transform -1 0 36432 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _548__223
timestamp 1666464484
transform -1 0 37536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _548_
timestamp 1666464484
transform 1 0 37260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _549_
timestamp 1666464484
transform -1 0 36432 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _549__224
timestamp 1666464484
transform -1 0 37444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _550_
timestamp 1666464484
transform 1 0 34500 0 -1 53312
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _550__225
timestamp 1666464484
transform 1 0 33764 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4140 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform -1 0 28520 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform -1 0 29900 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31740 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1666464484
transform 1 0 33764 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1666464484
transform -1 0 34040 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1666464484
transform 1 0 35880 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1666464484
transform 1 0 37260 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1666464484
transform 1 0 38640 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1666464484
transform 1 0 45448 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1666464484
transform 1 0 44988 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1666464484
transform 1 0 42780 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1666464484
transform 1 0 44712 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1666464484
transform -1 0 46000 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1666464484
transform 1 0 46920 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1666464484
transform 1 0 48300 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1666464484
transform 1 0 49680 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 51520 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 52532 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1666464484
transform 1 0 53912 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1666464484
transform 1 0 55292 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  macro_7_37
timestamp 1666464484
transform -1 0 50600 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_38
timestamp 1666464484
transform -1 0 51888 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_39
timestamp 1666464484
transform -1 0 53360 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_40
timestamp 1666464484
transform -1 0 54648 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_41
timestamp 1666464484
transform -1 0 56856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_42
timestamp 1666464484
transform -1 0 6808 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_43
timestamp 1666464484
transform -1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_44
timestamp 1666464484
transform 1 0 8924 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_45
timestamp 1666464484
transform 1 0 29624 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_46
timestamp 1666464484
transform -1 0 31648 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_47
timestamp 1666464484
transform -1 0 33948 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_48
timestamp 1666464484
transform -1 0 36432 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_49
timestamp 1666464484
transform -1 0 37536 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_50
timestamp 1666464484
transform -1 0 37536 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_51
timestamp 1666464484
transform -1 0 38824 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_52
timestamp 1666464484
transform 1 0 39284 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_53
timestamp 1666464484
transform -1 0 45816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_54
timestamp 1666464484
transform -1 0 47196 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_55
timestamp 1666464484
transform -1 0 46460 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_56
timestamp 1666464484
transform -1 0 47104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_57
timestamp 1666464484
transform -1 0 48484 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_58
timestamp 1666464484
transform -1 0 48576 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_59
timestamp 1666464484
transform -1 0 49956 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_60
timestamp 1666464484
transform -1 0 51244 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_61
timestamp 1666464484
transform -1 0 52716 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_62
timestamp 1666464484
transform -1 0 54004 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_63
timestamp 1666464484
transform -1 0 55476 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_64
timestamp 1666464484
transform -1 0 56488 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_65
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_66
timestamp 1666464484
transform 1 0 15824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_67
timestamp 1666464484
transform 1 0 17296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_68
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_69
timestamp 1666464484
transform -1 0 18768 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_70
timestamp 1666464484
transform 1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_71
timestamp 1666464484
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_72
timestamp 1666464484
transform 1 0 18584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_73
timestamp 1666464484
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_74
timestamp 1666464484
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_75
timestamp 1666464484
transform 1 0 19320 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_76
timestamp 1666464484
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_77
timestamp 1666464484
transform -1 0 20976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_78
timestamp 1666464484
transform 1 0 18676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_79
timestamp 1666464484
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_80
timestamp 1666464484
transform 1 0 17940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_81
timestamp 1666464484
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_82
timestamp 1666464484
transform 1 0 21344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_83
timestamp 1666464484
transform 1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_84
timestamp 1666464484
transform -1 0 22908 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_85
timestamp 1666464484
transform 1 0 19320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_86
timestamp 1666464484
transform 1 0 18584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_87
timestamp 1666464484
transform -1 0 23736 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_88
timestamp 1666464484
transform 1 0 19320 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_89
timestamp 1666464484
transform 1 0 22172 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_90
timestamp 1666464484
transform 1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_91
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_92
timestamp 1666464484
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_93
timestamp 1666464484
transform 1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_94
timestamp 1666464484
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_95
timestamp 1666464484
transform 1 0 21344 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_96
timestamp 1666464484
transform 1 0 22080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_97
timestamp 1666464484
transform -1 0 38916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_98
timestamp 1666464484
transform -1 0 39560 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_99
timestamp 1666464484
transform -1 0 40296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_100
timestamp 1666464484
transform -1 0 38180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_101
timestamp 1666464484
transform -1 0 38916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_102
timestamp 1666464484
transform -1 0 40296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_103
timestamp 1666464484
transform -1 0 39560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_104
timestamp 1666464484
transform -1 0 38088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_105
timestamp 1666464484
transform -1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_106
timestamp 1666464484
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_107
timestamp 1666464484
transform -1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_108
timestamp 1666464484
transform -1 0 40940 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_109
timestamp 1666464484
transform -1 0 39468 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_110
timestamp 1666464484
transform -1 0 40204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_111
timestamp 1666464484
transform -1 0 40848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_112
timestamp 1666464484
transform -1 0 40296 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_113
timestamp 1666464484
transform -1 0 42320 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_114
timestamp 1666464484
transform -1 0 41584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_115
timestamp 1666464484
transform -1 0 40940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_116
timestamp 1666464484
transform -1 0 42228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_117
timestamp 1666464484
transform -1 0 41676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_118
timestamp 1666464484
transform -1 0 43056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_119
timestamp 1666464484
transform -1 0 43056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_120
timestamp 1666464484
transform -1 0 42320 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_121
timestamp 1666464484
transform -1 0 43700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_122
timestamp 1666464484
transform -1 0 42964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_123
timestamp 1666464484
transform -1 0 43700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_124
timestamp 1666464484
transform -1 0 44436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_125
timestamp 1666464484
transform -1 0 43608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_126
timestamp 1666464484
transform -1 0 45080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_127
timestamp 1666464484
transform -1 0 44344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_128
timestamp 1666464484
transform -1 0 44436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_129
timestamp 1666464484
transform -1 0 44988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_130
timestamp 1666464484
transform -1 0 45816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_131
timestamp 1666464484
transform -1 0 46460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_132
timestamp 1666464484
transform -1 0 45816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_133
timestamp 1666464484
transform -1 0 45264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_134
timestamp 1666464484
transform -1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_135
timestamp 1666464484
transform -1 0 46460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_136
timestamp 1666464484
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_137
timestamp 1666464484
transform -1 0 47104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_138
timestamp 1666464484
transform -1 0 47196 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_139
timestamp 1666464484
transform -1 0 47748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_140
timestamp 1666464484
transform -1 0 48576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_141
timestamp 1666464484
transform -1 0 49220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_142
timestamp 1666464484
transform -1 0 48576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_143
timestamp 1666464484
transform -1 0 48024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_144
timestamp 1666464484
transform -1 0 49956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_145
timestamp 1666464484
transform -1 0 49220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_146
timestamp 1666464484
transform -1 0 50600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_147
timestamp 1666464484
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_148
timestamp 1666464484
transform -1 0 49956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_149
timestamp 1666464484
transform -1 0 50508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_150
timestamp 1666464484
transform -1 0 51336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_151
timestamp 1666464484
transform -1 0 51980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_152
timestamp 1666464484
transform -1 0 51336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_153
timestamp 1666464484
transform -1 0 50784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_154
timestamp 1666464484
transform -1 0 52716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_155
timestamp 1666464484
transform -1 0 51980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_156
timestamp 1666464484
transform -1 0 53360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_157
timestamp 1666464484
transform -1 0 52624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_158
timestamp 1666464484
transform -1 0 52716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_159
timestamp 1666464484
transform -1 0 53268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_160
timestamp 1666464484
transform -1 0 54096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_161
timestamp 1666464484
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_162
timestamp 1666464484
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_163
timestamp 1666464484
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_164
timestamp 1666464484
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_165
timestamp 1666464484
transform 1 0 8924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_166
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_167
timestamp 1666464484
transform 1 0 9752 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_168
timestamp 1666464484
transform -1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_169
timestamp 1666464484
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_170
timestamp 1666464484
transform 1 0 10396 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_171
timestamp 1666464484
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_172
timestamp 1666464484
transform 1 0 11040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_173
timestamp 1666464484
transform -1 0 11960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_174
timestamp 1666464484
transform 1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_175
timestamp 1666464484
transform -1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_176
timestamp 1666464484
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_177
timestamp 1666464484
transform 1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_178
timestamp 1666464484
transform -1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_179
timestamp 1666464484
transform 1 0 12420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_180
timestamp 1666464484
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_181
timestamp 1666464484
transform 1 0 13064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_182
timestamp 1666464484
transform -1 0 14444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_183
timestamp 1666464484
transform 1 0 13800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_184
timestamp 1666464484
transform 1 0 13800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_185
timestamp 1666464484
transform -1 0 15272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_186
timestamp 1666464484
transform 1 0 14444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_187
timestamp 1666464484
transform 1 0 14444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_188
timestamp 1666464484
transform -1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_189
timestamp 1666464484
transform 1 0 15272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_190
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_191
timestamp 1666464484
transform -1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_192
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_193
timestamp 1666464484
transform -1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_226
timestamp 1666464484
transform -1 0 4968 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_227
timestamp 1666464484
transform -1 0 6164 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_228
timestamp 1666464484
transform -1 0 7728 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_229
timestamp 1666464484
transform -1 0 9108 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_230
timestamp 1666464484
transform -1 0 10488 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_231
timestamp 1666464484
transform -1 0 11868 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_232
timestamp 1666464484
transform -1 0 13248 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_233
timestamp 1666464484
transform -1 0 14628 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_234
timestamp 1666464484
transform -1 0 16008 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_235
timestamp 1666464484
transform -1 0 17388 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_236
timestamp 1666464484
transform -1 0 18768 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_237
timestamp 1666464484
transform -1 0 20148 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_238
timestamp 1666464484
transform -1 0 21528 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_239
timestamp 1666464484
transform -1 0 22908 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_240
timestamp 1666464484
transform -1 0 24288 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_241
timestamp 1666464484
transform 1 0 24840 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_242
timestamp 1666464484
transform -1 0 27048 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_243
timestamp 1666464484
transform 1 0 26404 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_244
timestamp 1666464484
transform -1 0 30636 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_245
timestamp 1666464484
transform -1 0 31188 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_246
timestamp 1666464484
transform -1 0 35420 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_247
timestamp 1666464484
transform -1 0 35788 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_248
timestamp 1666464484
transform -1 0 35696 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_249
timestamp 1666464484
transform -1 0 37076 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_250
timestamp 1666464484
transform -1 0 38180 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_251
timestamp 1666464484
transform -1 0 43700 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_252
timestamp 1666464484
transform -1 0 45080 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_253
timestamp 1666464484
transform -1 0 46368 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_254
timestamp 1666464484
transform -1 0 43700 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_255
timestamp 1666464484
transform -1 0 45908 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_256
timestamp 1666464484
transform -1 0 47840 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_257
timestamp 1666464484
transform -1 0 47748 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_7_258
timestamp 1666464484
transform -1 0 49128 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1666464484
transform -1 0 5888 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1666464484
transform -1 0 18860 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1666464484
transform -1 0 20240 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1666464484
transform -1 0 21620 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1666464484
transform -1 0 23276 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1666464484
transform -1 0 23000 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1666464484
transform 1 0 25852 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1666464484
transform 1 0 30360 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1666464484
transform -1 0 29348 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1666464484
transform -1 0 10580 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1666464484
transform -1 0 11960 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1666464484
transform -1 0 13340 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1666464484
transform -1 0 14720 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1666464484
transform -1 0 16100 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1666464484
transform -1 0 17480 0 -1 57664
box -38 -48 406 592
<< labels >>
flabel metal2 s 3698 59200 3754 60000 0 FreeSans 224 90 0 0 io_active
port 0 nsew signal input
flabel metal2 s 4158 59200 4214 60000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 17958 59200 18014 60000 0 FreeSans 224 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s 19338 59200 19394 60000 0 FreeSans 224 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal2 s 20718 59200 20774 60000 0 FreeSans 224 90 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 22098 59200 22154 60000 0 FreeSans 224 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 23478 59200 23534 60000 0 FreeSans 224 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal2 s 24858 59200 24914 60000 0 FreeSans 224 90 0 0 io_in[15]
port 7 nsew signal input
flabel metal2 s 26238 59200 26294 60000 0 FreeSans 224 90 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 27618 59200 27674 60000 0 FreeSans 224 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 28998 59200 29054 60000 0 FreeSans 224 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 30378 59200 30434 60000 0 FreeSans 224 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal2 s 5538 59200 5594 60000 0 FreeSans 224 90 0 0 io_in[1]
port 12 nsew signal input
flabel metal2 s 31758 59200 31814 60000 0 FreeSans 224 90 0 0 io_in[20]
port 13 nsew signal input
flabel metal2 s 33138 59200 33194 60000 0 FreeSans 224 90 0 0 io_in[21]
port 14 nsew signal input
flabel metal2 s 34518 59200 34574 60000 0 FreeSans 224 90 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 35898 59200 35954 60000 0 FreeSans 224 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 37278 59200 37334 60000 0 FreeSans 224 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 38658 59200 38714 60000 0 FreeSans 224 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 40038 59200 40094 60000 0 FreeSans 224 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal2 s 41418 59200 41474 60000 0 FreeSans 224 90 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 42798 59200 42854 60000 0 FreeSans 224 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 44178 59200 44234 60000 0 FreeSans 224 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 6918 59200 6974 60000 0 FreeSans 224 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal2 s 45558 59200 45614 60000 0 FreeSans 224 90 0 0 io_in[30]
port 24 nsew signal input
flabel metal2 s 46938 59200 46994 60000 0 FreeSans 224 90 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 48318 59200 48374 60000 0 FreeSans 224 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal2 s 49698 59200 49754 60000 0 FreeSans 224 90 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 51078 59200 51134 60000 0 FreeSans 224 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 52458 59200 52514 60000 0 FreeSans 224 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal2 s 53838 59200 53894 60000 0 FreeSans 224 90 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 55218 59200 55274 60000 0 FreeSans 224 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 8298 59200 8354 60000 0 FreeSans 224 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal2 s 9678 59200 9734 60000 0 FreeSans 224 90 0 0 io_in[4]
port 33 nsew signal input
flabel metal2 s 11058 59200 11114 60000 0 FreeSans 224 90 0 0 io_in[5]
port 34 nsew signal input
flabel metal2 s 12438 59200 12494 60000 0 FreeSans 224 90 0 0 io_in[6]
port 35 nsew signal input
flabel metal2 s 13818 59200 13874 60000 0 FreeSans 224 90 0 0 io_in[7]
port 36 nsew signal input
flabel metal2 s 15198 59200 15254 60000 0 FreeSans 224 90 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 16578 59200 16634 60000 0 FreeSans 224 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 4618 59200 4674 60000 0 FreeSans 224 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal2 s 18418 59200 18474 60000 0 FreeSans 224 90 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal2 s 19798 59200 19854 60000 0 FreeSans 224 90 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal2 s 21178 59200 21234 60000 0 FreeSans 224 90 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal2 s 22558 59200 22614 60000 0 FreeSans 224 90 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal2 s 23938 59200 23994 60000 0 FreeSans 224 90 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 25318 59200 25374 60000 0 FreeSans 224 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal2 s 26698 59200 26754 60000 0 FreeSans 224 90 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 28078 59200 28134 60000 0 FreeSans 224 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 29458 59200 29514 60000 0 FreeSans 224 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 30838 59200 30894 60000 0 FreeSans 224 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal2 s 5998 59200 6054 60000 0 FreeSans 224 90 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal2 s 32218 59200 32274 60000 0 FreeSans 224 90 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal2 s 33598 59200 33654 60000 0 FreeSans 224 90 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 34978 59200 35034 60000 0 FreeSans 224 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 36358 59200 36414 60000 0 FreeSans 224 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 37738 59200 37794 60000 0 FreeSans 224 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal2 s 39118 59200 39174 60000 0 FreeSans 224 90 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal2 s 40498 59200 40554 60000 0 FreeSans 224 90 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 41878 59200 41934 60000 0 FreeSans 224 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal2 s 43258 59200 43314 60000 0 FreeSans 224 90 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal2 s 44638 59200 44694 60000 0 FreeSans 224 90 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 7378 59200 7434 60000 0 FreeSans 224 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal2 s 46018 59200 46074 60000 0 FreeSans 224 90 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal2 s 47398 59200 47454 60000 0 FreeSans 224 90 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal2 s 48778 59200 48834 60000 0 FreeSans 224 90 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal2 s 50158 59200 50214 60000 0 FreeSans 224 90 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal2 s 51538 59200 51594 60000 0 FreeSans 224 90 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal2 s 52918 59200 52974 60000 0 FreeSans 224 90 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal2 s 54298 59200 54354 60000 0 FreeSans 224 90 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal2 s 55678 59200 55734 60000 0 FreeSans 224 90 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 8758 59200 8814 60000 0 FreeSans 224 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal2 s 10138 59200 10194 60000 0 FreeSans 224 90 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal2 s 11518 59200 11574 60000 0 FreeSans 224 90 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal2 s 12898 59200 12954 60000 0 FreeSans 224 90 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 14278 59200 14334 60000 0 FreeSans 224 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 15658 59200 15714 60000 0 FreeSans 224 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 17038 59200 17094 60000 0 FreeSans 224 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal2 s 5078 59200 5134 60000 0 FreeSans 224 90 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal2 s 18878 59200 18934 60000 0 FreeSans 224 90 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal2 s 20258 59200 20314 60000 0 FreeSans 224 90 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal2 s 21638 59200 21694 60000 0 FreeSans 224 90 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal2 s 23018 59200 23074 60000 0 FreeSans 224 90 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal2 s 24398 59200 24454 60000 0 FreeSans 224 90 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal2 s 25778 59200 25834 60000 0 FreeSans 224 90 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal2 s 27158 59200 27214 60000 0 FreeSans 224 90 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 28538 59200 28594 60000 0 FreeSans 224 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal2 s 29918 59200 29974 60000 0 FreeSans 224 90 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal2 s 31298 59200 31354 60000 0 FreeSans 224 90 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 6458 59200 6514 60000 0 FreeSans 224 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 32678 59200 32734 60000 0 FreeSans 224 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal2 s 34058 59200 34114 60000 0 FreeSans 224 90 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 35438 59200 35494 60000 0 FreeSans 224 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal2 s 36818 59200 36874 60000 0 FreeSans 224 90 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 38198 59200 38254 60000 0 FreeSans 224 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 39578 59200 39634 60000 0 FreeSans 224 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal2 s 40958 59200 41014 60000 0 FreeSans 224 90 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 42338 59200 42394 60000 0 FreeSans 224 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 43718 59200 43774 60000 0 FreeSans 224 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal2 s 45098 59200 45154 60000 0 FreeSans 224 90 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 7838 59200 7894 60000 0 FreeSans 224 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal2 s 46478 59200 46534 60000 0 FreeSans 224 90 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal2 s 47858 59200 47914 60000 0 FreeSans 224 90 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal2 s 49238 59200 49294 60000 0 FreeSans 224 90 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal2 s 50618 59200 50674 60000 0 FreeSans 224 90 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal2 s 51998 59200 52054 60000 0 FreeSans 224 90 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal2 s 53378 59200 53434 60000 0 FreeSans 224 90 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 54758 59200 54814 60000 0 FreeSans 224 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal2 s 56138 59200 56194 60000 0 FreeSans 224 90 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal2 s 9218 59200 9274 60000 0 FreeSans 224 90 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal2 s 10598 59200 10654 60000 0 FreeSans 224 90 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 11978 59200 12034 60000 0 FreeSans 224 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 13358 59200 13414 60000 0 FreeSans 224 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal2 s 14738 59200 14794 60000 0 FreeSans 224 90 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 16118 59200 16174 60000 0 FreeSans 224 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal2 s 17498 59200 17554 60000 0 FreeSans 224 90 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 115 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 116 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 117 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 118 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 119 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 120 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 121 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 122 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 123 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 124 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 125 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 126 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 127 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 128 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 129 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 130 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 131 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 132 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 133 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 134 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 135 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 136 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 137 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 138 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 139 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 140 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 141 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 142 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 143 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 144 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 145 nsew signal input
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 146 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 147 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 148 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 149 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 150 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 151 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 152 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 153 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 154 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 155 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 156 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 157 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 158 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 159 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 160 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 161 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 162 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 163 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 164 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 165 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 166 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 167 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 168 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 169 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 170 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 171 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 172 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 173 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 174 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 175 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 176 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 177 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 178 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 179 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 180 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 181 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 182 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 183 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 184 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 185 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 186 nsew signal input
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 187 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 188 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 189 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 190 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 191 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 192 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 193 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 194 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 195 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 196 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 197 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 198 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 199 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 200 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 201 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 202 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 203 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 204 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 205 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 206 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 207 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 208 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 209 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 210 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 211 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 212 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 213 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 214 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 215 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 216 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 217 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 218 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 219 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 220 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 221 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 222 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 223 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 224 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 225 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 226 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 227 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 228 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 229 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 230 nsew signal input
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 231 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 232 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 233 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 234 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 235 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 236 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 237 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 238 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 239 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 240 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 241 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 242 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 243 nsew signal tristate
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 244 nsew signal tristate
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 245 nsew signal tristate
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 246 nsew signal tristate
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 247 nsew signal tristate
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 248 nsew signal tristate
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 249 nsew signal tristate
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 250 nsew signal tristate
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 251 nsew signal tristate
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 252 nsew signal tristate
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 253 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 254 nsew signal tristate
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 255 nsew signal tristate
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 256 nsew signal tristate
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 257 nsew signal tristate
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 258 nsew signal tristate
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 259 nsew signal tristate
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 260 nsew signal tristate
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 261 nsew signal tristate
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 262 nsew signal tristate
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 263 nsew signal tristate
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 264 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 265 nsew signal tristate
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 266 nsew signal tristate
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 267 nsew signal tristate
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 268 nsew signal tristate
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 269 nsew signal tristate
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 270 nsew signal tristate
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 271 nsew signal tristate
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 272 nsew signal tristate
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 273 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 274 nsew signal tristate
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 275 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 276 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 277 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 278 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 279 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 280 nsew signal tristate
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 281 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 282 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 283 nsew signal tristate
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 284 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 285 nsew signal tristate
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 286 nsew signal tristate
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 287 nsew signal tristate
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 288 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 289 nsew signal tristate
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 290 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 291 nsew signal tristate
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 292 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 293 nsew signal tristate
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 294 nsew signal tristate
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 295 nsew signal tristate
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 296 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 297 nsew signal tristate
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 298 nsew signal tristate
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 299 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 300 nsew signal tristate
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 301 nsew signal tristate
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 302 nsew signal tristate
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 303 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 304 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 305 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 306 nsew signal tristate
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 307 nsew signal tristate
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 308 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 309 nsew signal tristate
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 310 nsew signal tristate
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 311 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 312 nsew signal tristate
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 313 nsew signal tristate
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 314 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 315 nsew signal tristate
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 316 nsew signal tristate
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 317 nsew signal tristate
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 318 nsew signal tristate
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 319 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 320 nsew signal tristate
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 321 nsew signal tristate
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 322 nsew signal tristate
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 323 nsew signal tristate
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 324 nsew signal tristate
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 325 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 326 nsew signal tristate
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 327 nsew signal tristate
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 328 nsew signal tristate
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 329 nsew signal tristate
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 330 nsew signal tristate
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 331 nsew signal tristate
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 332 nsew signal tristate
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 333 nsew signal tristate
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 334 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 335 nsew signal tristate
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 336 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 337 nsew signal tristate
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 338 nsew signal tristate
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 339 nsew signal tristate
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 340 nsew signal tristate
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 341 nsew signal tristate
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 342 nsew signal tristate
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 343 nsew signal tristate
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 344 nsew signal tristate
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 345 nsew signal tristate
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 346 nsew signal tristate
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 347 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 348 nsew signal tristate
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 349 nsew signal tristate
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 350 nsew signal tristate
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 351 nsew signal tristate
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 352 nsew signal tristate
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 353 nsew signal tristate
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 354 nsew signal tristate
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 355 nsew signal tristate
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 356 nsew signal tristate
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 357 nsew signal tristate
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 358 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 359 nsew signal tristate
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 360 nsew signal tristate
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 361 nsew signal tristate
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 362 nsew signal tristate
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 363 nsew signal tristate
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 364 nsew signal tristate
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 365 nsew signal tristate
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 366 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 367 nsew signal tristate
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 368 nsew signal tristate
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 369 nsew signal tristate
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 370 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 371 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 372 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 373 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 374 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 375 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 376 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 377 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 378 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 379 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 380 nsew signal input
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 381 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 382 nsew signal input
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 383 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 384 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 385 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 386 nsew signal input
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 387 nsew signal input
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 388 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 389 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 390 nsew signal input
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 391 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 392 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 393 nsew signal input
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 394 nsew signal input
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 395 nsew signal input
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 396 nsew signal input
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 397 nsew signal input
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 398 nsew signal input
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 399 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 400 nsew signal input
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 401 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 402 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 403 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 404 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 405 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 406 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 407 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 408 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 409 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 410 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 411 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 412 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 413 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 414 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 415 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 416 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 417 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 418 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 419 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 420 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 421 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 422 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 423 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 424 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 425 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 426 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 427 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 428 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 429 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 430 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 431 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 432 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 433 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 434 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 435 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 436 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 437 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 438 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 439 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 440 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 441 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 442 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 443 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 444 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 445 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 446 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 447 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 448 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 449 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 450 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 451 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 452 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 453 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 454 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 455 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 456 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 457 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 458 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 459 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 460 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 461 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 462 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 463 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 464 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 465 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 466 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 467 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 468 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 469 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 470 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 471 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 472 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 473 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 474 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 475 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 476 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 477 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 478 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 479 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 480 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 481 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 482 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 483 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 484 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 485 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 486 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 487 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 488 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 489 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 490 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 491 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 492 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 493 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 494 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 495 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 496 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 497 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 498 nsew signal input
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 500 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 500 nsew ground bidirectional
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wb_clk_i
port 501 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wb_rst_i
port 502 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 503 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 504 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 505 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 506 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 507 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 508 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 509 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 510 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 511 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 512 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 513 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 514 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 515 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 516 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 517 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 518 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 519 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 520 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 521 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 522 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 523 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 524 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 525 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 526 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 527 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 528 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 529 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 530 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 531 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 532 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 533 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 534 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 535 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 536 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 537 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 538 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 539 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 540 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 541 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 542 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 543 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 544 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 545 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 546 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 547 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 548 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 549 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 550 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 551 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 552 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 553 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 554 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 555 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 556 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 557 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 558 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 559 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 560 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 561 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 562 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 563 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 564 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 565 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 566 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 567 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 568 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 569 nsew signal tristate
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 570 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 571 nsew signal tristate
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 572 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 573 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 574 nsew signal tristate
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 575 nsew signal tristate
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 576 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 577 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 578 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 579 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 580 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 581 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 582 nsew signal tristate
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 583 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 584 nsew signal tristate
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 585 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 586 nsew signal tristate
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 587 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 588 nsew signal tristate
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 589 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 590 nsew signal tristate
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 591 nsew signal tristate
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 592 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 593 nsew signal tristate
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 594 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 595 nsew signal tristate
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 596 nsew signal tristate
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 597 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 598 nsew signal tristate
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 599 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 600 nsew signal tristate
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 601 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 602 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 603 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 604 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 605 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_we_i
port 606 nsew signal input
rlabel metal1 29992 57120 29992 57120 0 vccd1
rlabel metal1 29992 57664 29992 57664 0 vssd1
rlabel metal2 36202 55114 36202 55114 0 _000_
rlabel metal2 34638 56066 34638 56066 0 _001_
rlabel metal1 30268 56338 30268 56338 0 _002_
rlabel metal1 27370 55590 27370 55590 0 _003_
rlabel metal1 35788 54706 35788 54706 0 _004_
rlabel metal1 33281 54842 33281 54842 0 _005_
rlabel metal1 29302 54298 29302 54298 0 _006_
rlabel metal1 33902 54230 33902 54230 0 _007_
rlabel metal2 33350 54332 33350 54332 0 _008_
rlabel metal1 33028 54298 33028 54298 0 _009_
rlabel metal2 32338 54876 32338 54876 0 _010_
rlabel metal1 33304 53686 33304 53686 0 _011_
rlabel metal1 29256 55250 29256 55250 0 _012_
rlabel metal1 30130 55352 30130 55352 0 _013_
rlabel metal2 30038 54774 30038 54774 0 _014_
rlabel metal1 28336 55726 28336 55726 0 _015_
rlabel metal2 33994 55998 33994 55998 0 _016_
rlabel metal2 28290 56100 28290 56100 0 _017_
rlabel metal1 28198 56406 28198 56406 0 _018_
rlabel metal1 28152 56474 28152 56474 0 _019_
rlabel metal2 44390 56134 44390 56134 0 _020_
rlabel metal1 43056 56270 43056 56270 0 _021_
rlabel metal2 37030 55845 37030 55845 0 _022_
rlabel metal1 38272 56202 38272 56202 0 _023_
rlabel metal1 43562 55182 43562 55182 0 _024_
rlabel metal1 39146 55148 39146 55148 0 _025_
rlabel metal2 38962 55658 38962 55658 0 _026_
rlabel metal1 42090 55590 42090 55590 0 _027_
rlabel metal2 42274 54672 42274 54672 0 _028_
rlabel metal2 41446 55080 41446 55080 0 _029_
rlabel metal2 40802 54842 40802 54842 0 _030_
rlabel metal1 40756 53958 40756 53958 0 _031_
rlabel metal1 39054 55760 39054 55760 0 _032_
rlabel metal1 38686 56270 38686 56270 0 _033_
rlabel metal1 37858 55692 37858 55692 0 _034_
rlabel metal1 39054 56338 39054 56338 0 _035_
rlabel metal1 39652 56338 39652 56338 0 _036_
rlabel metal1 36570 56236 36570 56236 0 _037_
rlabel metal1 37306 56406 37306 56406 0 _038_
rlabel metal1 36294 56474 36294 56474 0 _039_
rlabel metal2 34454 56372 34454 56372 0 _040_
rlabel metal1 31878 56338 31878 56338 0 _041_
rlabel metal1 31832 56474 31832 56474 0 _042_
rlabel metal1 24731 56814 24731 56814 0 _043_
rlabel metal1 37122 56678 37122 56678 0 _044_
rlabel metal2 40342 56202 40342 56202 0 _045_
rlabel metal2 40526 56644 40526 56644 0 _046_
rlabel metal1 40020 57562 40020 57562 0 _047_
rlabel metal2 24058 56610 24058 56610 0 _048_
rlabel metal2 24334 56576 24334 56576 0 _049_
rlabel metal1 32522 54638 32522 54638 0 _050_
rlabel metal1 32844 54774 32844 54774 0 _051_
rlabel metal2 33810 57120 33810 57120 0 _052_
rlabel metal1 33074 56338 33074 56338 0 _053_
rlabel metal2 32706 56746 32706 56746 0 _054_
rlabel metal2 41354 54468 41354 54468 0 _055_
rlabel metal1 41814 54842 41814 54842 0 _056_
rlabel metal1 42320 56814 42320 56814 0 _057_
rlabel viali 41430 56338 41430 56338 0 _058_
rlabel metal2 41170 55981 41170 55981 0 _059_
rlabel metal2 25714 55692 25714 55692 0 _060_
rlabel metal2 25622 55930 25622 55930 0 _061_
rlabel metal1 31602 55658 31602 55658 0 _062_
rlabel metal1 32637 55794 32637 55794 0 _063_
rlabel metal1 30636 55318 30636 55318 0 _064_
rlabel metal1 30912 55386 30912 55386 0 _065_
rlabel via1 30310 55386 30310 55386 0 _066_
rlabel metal2 27370 55862 27370 55862 0 _067_
rlabel metal1 40618 56406 40618 56406 0 _068_
rlabel metal2 40986 56134 40986 56134 0 _069_
rlabel metal2 39698 54842 39698 54842 0 _070_
rlabel metal1 40020 54842 40020 54842 0 _071_
rlabel metal2 40066 55148 40066 55148 0 _072_
rlabel via2 40710 56219 40710 56219 0 _073_
rlabel metal2 27094 55930 27094 55930 0 _074_
rlabel metal1 25254 55760 25254 55760 0 _075_
rlabel metal1 28934 54638 28934 54638 0 _076_
rlabel metal2 28750 54876 28750 54876 0 _077_
rlabel metal1 29348 54774 29348 54774 0 _078_
rlabel metal1 30866 54230 30866 54230 0 _079_
rlabel metal2 28474 55828 28474 55828 0 _080_
rlabel metal2 28566 55692 28566 55692 0 _081_
rlabel metal1 28750 54842 28750 54842 0 _082_
rlabel metal2 37674 56032 37674 56032 0 _083_
rlabel metal1 38042 56270 38042 56270 0 _084_
rlabel metal2 37306 56644 37306 56644 0 _085_
rlabel metal2 44206 57052 44206 57052 0 _086_
rlabel metal1 37536 56814 37536 56814 0 _087_
rlabel metal2 37398 56695 37398 56695 0 _088_
rlabel metal2 21942 57324 21942 57324 0 _089_
rlabel metal1 37030 2414 37030 2414 0 _090_
rlabel metal1 28980 2414 28980 2414 0 _091_
rlabel metal2 26266 7072 26266 7072 0 _092_
rlabel metal2 25438 5372 25438 5372 0 _093_
rlabel metal2 22678 4012 22678 4012 0 _094_
rlabel metal1 22862 2856 22862 2856 0 _095_
rlabel metal2 22218 3570 22218 3570 0 _096_
rlabel metal2 24058 4318 24058 4318 0 _097_
rlabel metal2 26818 6494 26818 6494 0 _098_
rlabel metal1 27140 5270 27140 5270 0 _099_
rlabel metal2 27830 4828 27830 4828 0 _100_
rlabel metal1 28198 3604 28198 3604 0 _101_
rlabel metal1 24012 3910 24012 3910 0 _102_
rlabel metal1 24518 2550 24518 2550 0 _103_
rlabel metal1 25760 2482 25760 2482 0 _104_
rlabel metal1 26588 2550 26588 2550 0 _105_
rlabel metal1 29486 4046 29486 4046 0 _106_
rlabel metal2 29486 6766 29486 6766 0 _107_
rlabel metal1 29900 5270 29900 5270 0 _108_
rlabel metal1 29532 2346 29532 2346 0 _109_
rlabel metal1 30084 2618 30084 2618 0 _110_
rlabel metal1 28658 2550 28658 2550 0 _111_
rlabel metal2 33442 5950 33442 5950 0 _112_
rlabel metal2 30958 6460 30958 6460 0 _113_
rlabel metal1 33350 2618 33350 2618 0 _114_
rlabel metal1 33626 3434 33626 3434 0 _115_
rlabel metal1 35006 2618 35006 2618 0 _116_
rlabel metal2 32338 5610 32338 5610 0 _117_
rlabel metal1 33350 4692 33350 4692 0 _118_
rlabel metal2 34822 5916 34822 5916 0 _119_
rlabel metal1 36064 2618 36064 2618 0 _120_
rlabel metal2 36202 4318 36202 4318 0 _121_
rlabel metal1 37444 2618 37444 2618 0 _122_
rlabel metal1 37996 2618 37996 2618 0 _123_
rlabel metal1 35282 56372 35282 56372 0 _124_
rlabel metal1 3680 57562 3680 57562 0 io_active
rlabel metal1 28612 54162 28612 54162 0 io_in[18]
rlabel metal1 30084 57562 30084 57562 0 io_in[19]
rlabel metal2 31786 58320 31786 58320 0 io_in[20]
rlabel metal1 33764 54162 33764 54162 0 io_in[21]
rlabel metal1 33902 56440 33902 56440 0 io_in[22]
rlabel metal2 35926 55522 35926 55522 0 io_in[23]
rlabel metal1 37398 57358 37398 57358 0 io_in[24]
rlabel metal1 39284 57426 39284 57426 0 io_in[25]
rlabel metal2 45678 56865 45678 56865 0 io_in[26]
rlabel metal1 45218 55760 45218 55760 0 io_in[27]
rlabel metal2 42826 58587 42826 58587 0 io_in[28]
rlabel metal1 44942 55284 44942 55284 0 io_in[29]
rlabel metal1 45724 57494 45724 57494 0 io_in[30]
rlabel metal2 46966 58320 46966 58320 0 io_in[31]
rlabel metal2 48346 58320 48346 58320 0 io_in[32]
rlabel metal2 49726 58320 49726 58320 0 io_in[33]
rlabel metal1 51290 57426 51290 57426 0 io_in[34]
rlabel via1 52578 57494 52578 57494 0 io_in[35]
rlabel metal1 53912 57426 53912 57426 0 io_in[36]
rlabel metal1 55292 57426 55292 57426 0 io_in[37]
rlabel metal1 5612 57562 5612 57562 0 io_out[0]
rlabel metal1 18768 57562 18768 57562 0 io_out[10]
rlabel metal1 20148 57562 20148 57562 0 io_out[11]
rlabel metal1 21482 57562 21482 57562 0 io_out[12]
rlabel metal2 23046 58116 23046 58116 0 io_out[13]
rlabel metal1 23598 57562 23598 57562 0 io_out[14]
rlabel metal1 25944 55930 25944 55930 0 io_out[15]
rlabel metal1 30590 57528 30590 57528 0 io_out[16]
rlabel metal1 29072 57562 29072 57562 0 io_out[17]
rlabel metal1 10488 57562 10488 57562 0 io_out[4]
rlabel metal1 11868 57562 11868 57562 0 io_out[5]
rlabel metal1 13248 57562 13248 57562 0 io_out[6]
rlabel metal1 14628 57562 14628 57562 0 io_out[7]
rlabel metal1 16008 57562 16008 57562 0 io_out[8]
rlabel metal1 17388 57562 17388 57562 0 io_out[9]
rlabel metal2 26174 1761 26174 1761 0 la_data_out[32]
rlabel metal1 25392 3366 25392 3366 0 la_data_out[33]
rlabel metal2 26726 3254 26726 3254 0 la_data_out[34]
rlabel metal1 26358 3910 26358 3910 0 la_data_out[35]
rlabel metal1 26496 3094 26496 3094 0 la_data_out[36]
rlabel metal2 27554 3492 27554 3492 0 la_data_out[37]
rlabel metal2 27830 1690 27830 1690 0 la_data_out[38]
rlabel metal2 28106 1520 28106 1520 0 la_data_out[39]
rlabel metal1 28428 3570 28428 3570 0 la_data_out[40]
rlabel metal2 28658 3254 28658 3254 0 la_data_out[41]
rlabel metal1 28014 3434 28014 3434 0 la_data_out[42]
rlabel metal1 29210 4012 29210 4012 0 la_data_out[43]
rlabel metal1 28980 2890 28980 2890 0 la_data_out[44]
rlabel metal2 29762 2404 29762 2404 0 la_data_out[45]
rlabel metal2 30038 3492 30038 3492 0 la_data_out[46]
rlabel metal2 30360 4692 30360 4692 0 la_data_out[47]
rlabel metal2 30590 1503 30590 1503 0 la_data_out[48]
rlabel metal1 30958 3570 30958 3570 0 la_data_out[49]
rlabel metal2 31142 1860 31142 1860 0 la_data_out[50]
rlabel metal2 31786 3978 31786 3978 0 la_data_out[51]
rlabel metal2 31694 3254 31694 3254 0 la_data_out[52]
rlabel metal2 31970 1860 31970 1860 0 la_data_out[53]
rlabel metal1 32936 3570 32936 3570 0 la_data_out[54]
rlabel metal1 33764 2890 33764 2890 0 la_data_out[55]
rlabel metal2 32798 2404 32798 2404 0 la_data_out[56]
rlabel metal1 33350 3162 33350 3162 0 la_data_out[57]
rlabel metal2 33350 3254 33350 3254 0 la_data_out[58]
rlabel metal2 33626 1299 33626 1299 0 la_data_out[59]
rlabel metal2 33902 1435 33902 1435 0 la_data_out[60]
rlabel metal1 35052 3094 35052 3094 0 la_data_out[61]
rlabel metal2 34500 4012 34500 4012 0 la_data_out[62]
rlabel metal2 34730 1639 34730 1639 0 la_data_out[63]
rlabel metal2 11086 57086 11086 57086 0 net1
rlabel metal1 40526 56678 40526 56678 0 net10
rlabel metal1 36892 4046 36892 4046 0 net100
rlabel metal2 36110 1299 36110 1299 0 net101
rlabel metal1 37812 3094 37812 3094 0 net102
rlabel metal1 36984 3434 36984 3434 0 net103
rlabel metal1 37398 3706 37398 3706 0 net104
rlabel metal2 37214 1622 37214 1622 0 net105
rlabel metal2 37490 1367 37490 1367 0 net106
rlabel metal2 37766 1554 37766 1554 0 net107
rlabel metal1 39376 2890 39376 2890 0 net108
rlabel metal1 38778 3910 38778 3910 0 net109
rlabel metal2 42734 56474 42734 56474 0 net11
rlabel metal1 39284 3570 39284 3570 0 net110
rlabel metal1 39744 3434 39744 3434 0 net111
rlabel metal1 39606 4046 39606 4046 0 net112
rlabel metal2 39422 1656 39422 1656 0 net113
rlabel metal1 40526 3026 40526 3026 0 net114
rlabel metal1 40342 3978 40342 3978 0 net115
rlabel metal2 40250 1860 40250 1860 0 net116
rlabel metal2 40526 2200 40526 2200 0 net117
rlabel metal2 40802 1554 40802 1554 0 net118
rlabel metal1 42113 2822 42113 2822 0 net119
rlabel metal1 39054 55284 39054 55284 0 net12
rlabel metal2 41354 2166 41354 2166 0 net120
rlabel metal2 41630 1622 41630 1622 0 net121
rlabel metal2 41906 2098 41906 2098 0 net122
rlabel metal2 42182 1860 42182 1860 0 net123
rlabel metal2 42458 1656 42458 1656 0 net124
rlabel metal2 42734 2200 42734 2200 0 net125
rlabel metal2 43010 1588 43010 1588 0 net126
rlabel metal2 43286 1826 43286 1826 0 net127
rlabel metal2 43562 2132 43562 2132 0 net128
rlabel metal2 43838 1792 43838 1792 0 net129
rlabel metal1 37996 54638 37996 54638 0 net13
rlabel metal2 44114 1622 44114 1622 0 net130
rlabel metal2 44390 1554 44390 1554 0 net131
rlabel metal2 44666 1860 44666 1860 0 net132
rlabel metal2 44942 2132 44942 2132 0 net133
rlabel metal2 45218 1656 45218 1656 0 net134
rlabel metal2 45494 1826 45494 1826 0 net135
rlabel metal2 45770 1554 45770 1554 0 net136
rlabel metal2 46046 1792 46046 1792 0 net137
rlabel metal2 46322 2132 46322 2132 0 net138
rlabel metal2 46598 1826 46598 1826 0 net139
rlabel metal2 44114 56304 44114 56304 0 net14
rlabel metal2 46874 1622 46874 1622 0 net140
rlabel metal2 47150 1690 47150 1690 0 net141
rlabel metal2 47426 1792 47426 1792 0 net142
rlabel metal2 47702 2132 47702 2132 0 net143
rlabel metal2 47978 1656 47978 1656 0 net144
rlabel metal2 48254 1826 48254 1826 0 net145
rlabel metal2 48530 1588 48530 1588 0 net146
rlabel metal2 48806 1792 48806 1792 0 net147
rlabel metal2 49082 2132 49082 2132 0 net148
rlabel metal2 49358 1826 49358 1826 0 net149
rlabel metal1 44574 56202 44574 56202 0 net15
rlabel metal2 49634 1622 49634 1622 0 net150
rlabel metal2 49910 1690 49910 1690 0 net151
rlabel metal2 50186 1792 50186 1792 0 net152
rlabel metal2 50462 1299 50462 1299 0 net153
rlabel metal2 50738 1554 50738 1554 0 net154
rlabel metal2 51014 1826 51014 1826 0 net155
rlabel metal2 51290 1656 51290 1656 0 net156
rlabel metal2 51566 1792 51566 1792 0 net157
rlabel metal2 51842 2132 51842 2132 0 net158
rlabel metal2 52118 1826 52118 1826 0 net159
rlabel metal2 44022 56950 44022 56950 0 net16
rlabel metal2 52394 1622 52394 1622 0 net160
rlabel metal2 7682 1588 7682 1588 0 net161
rlabel metal2 8234 1588 8234 1588 0 net162
rlabel metal2 8602 1792 8602 1792 0 net163
rlabel metal2 8970 1588 8970 1588 0 net164
rlabel metal2 9338 1792 9338 1792 0 net165
rlabel metal2 9706 1588 9706 1588 0 net166
rlabel metal2 9982 1792 9982 1792 0 net167
rlabel metal2 10258 2132 10258 2132 0 net168
rlabel metal2 10534 1656 10534 1656 0 net169
rlabel metal1 45126 57358 45126 57358 0 net17
rlabel metal2 10810 1792 10810 1792 0 net170
rlabel metal2 11086 1588 11086 1588 0 net171
rlabel metal2 11362 1792 11362 1792 0 net172
rlabel metal2 11638 1792 11638 1792 0 net173
rlabel metal2 11914 1656 11914 1656 0 net174
rlabel metal2 12190 2132 12190 2132 0 net175
rlabel metal2 12466 1588 12466 1588 0 net176
rlabel metal2 12742 1792 12742 1792 0 net177
rlabel metal2 13018 2132 13018 2132 0 net178
rlabel metal2 13294 1656 13294 1656 0 net179
rlabel metal2 51290 57698 51290 57698 0 net18
rlabel metal2 13570 1792 13570 1792 0 net180
rlabel metal2 13846 1588 13846 1588 0 net181
rlabel metal2 14122 2132 14122 2132 0 net182
rlabel metal2 14398 1792 14398 1792 0 net183
rlabel metal2 14674 1656 14674 1656 0 net184
rlabel metal2 14950 2132 14950 2132 0 net185
rlabel metal2 15226 1792 15226 1792 0 net186
rlabel metal2 15502 1588 15502 1588 0 net187
rlabel metal2 15778 2132 15778 2132 0 net188
rlabel metal2 16054 1792 16054 1792 0 net189
rlabel metal2 51106 56542 51106 56542 0 net19
rlabel metal2 16330 1792 16330 1792 0 net190
rlabel metal2 16606 2132 16606 2132 0 net191
rlabel metal2 16882 1622 16882 1622 0 net192
rlabel metal2 17158 2336 17158 2336 0 net193
rlabel metal2 25254 5712 25254 5712 0 net194
rlabel metal2 22494 3740 22494 3740 0 net195
rlabel metal2 22126 3842 22126 3842 0 net196
rlabel metal1 23414 2618 23414 2618 0 net197
rlabel metal2 22402 3264 22402 3264 0 net198
rlabel metal1 24518 5134 24518 5134 0 net199
rlabel metal1 31924 55046 31924 55046 0 net2
rlabel metal2 54142 57086 54142 57086 0 net20
rlabel metal2 26634 5984 26634 5984 0 net200
rlabel metal2 27646 5712 27646 5712 0 net201
rlabel metal2 28014 5372 28014 5372 0 net202
rlabel metal1 25438 2822 25438 2822 0 net203
rlabel metal1 25162 3570 25162 3570 0 net204
rlabel metal1 24840 2618 24840 2618 0 net205
rlabel metal1 26174 2618 26174 2618 0 net206
rlabel metal1 29118 4114 29118 4114 0 net207
rlabel metal2 29302 6528 29302 6528 0 net208
rlabel metal2 29394 5984 29394 5984 0 net209
rlabel metal2 50094 56542 50094 56542 0 net21
rlabel metal1 29854 2482 29854 2482 0 net210
rlabel metal1 30636 2618 30636 2618 0 net211
rlabel metal1 27830 2618 27830 2618 0 net212
rlabel metal2 33626 5678 33626 5678 0 net213
rlabel metal2 31786 6290 31786 6290 0 net214
rlabel metal1 32798 2550 32798 2550 0 net215
rlabel metal1 32890 2618 32890 2618 0 net216
rlabel metal2 34546 2788 34546 2788 0 net217
rlabel metal2 32154 5100 32154 5100 0 net218
rlabel metal2 33166 5712 33166 5712 0 net219
rlabel via2 6394 57443 6394 57443 0 net22
rlabel metal1 35006 5780 35006 5780 0 net220
rlabel metal1 36248 2550 36248 2550 0 net221
rlabel metal2 36386 4352 36386 4352 0 net222
rlabel metal2 37306 3468 37306 3468 0 net223
rlabel metal2 37214 4964 37214 4964 0 net224
rlabel metal1 34270 53006 34270 53006 0 net225
rlabel metal1 4692 57018 4692 57018 0 net226
rlabel metal1 5980 57018 5980 57018 0 net227
rlabel metal1 7452 57426 7452 57426 0 net228
rlabel metal1 8832 57018 8832 57018 0 net229
rlabel metal1 18814 57392 18814 57392 0 net23
rlabel metal1 10212 57018 10212 57018 0 net230
rlabel metal1 11592 57018 11592 57018 0 net231
rlabel metal1 12972 57018 12972 57018 0 net232
rlabel metal1 14352 57018 14352 57018 0 net233
rlabel metal1 15732 57018 15732 57018 0 net234
rlabel metal1 17112 57018 17112 57018 0 net235
rlabel metal1 18492 57018 18492 57018 0 net236
rlabel metal1 19964 57018 19964 57018 0 net237
rlabel metal1 21252 57018 21252 57018 0 net238
rlabel metal1 22632 56338 22632 56338 0 net239
rlabel metal2 20194 57664 20194 57664 0 net24
rlabel metal1 24012 55182 24012 55182 0 net240
rlabel metal1 25208 55182 25208 55182 0 net241
rlabel metal1 26772 54162 26772 54162 0 net242
rlabel metal1 27232 55182 27232 55182 0 net243
rlabel metal1 30084 53754 30084 53754 0 net244
rlabel metal1 30912 56338 30912 56338 0 net245
rlabel metal1 34776 56882 34776 56882 0 net246
rlabel metal1 35098 55182 35098 55182 0 net247
rlabel metal1 35420 54162 35420 54162 0 net248
rlabel metal1 36616 54842 36616 54842 0 net249
rlabel metal2 21850 57630 21850 57630 0 net25
rlabel metal1 37858 54162 37858 54162 0 net250
rlabel metal2 43470 57358 43470 57358 0 net251
rlabel metal2 44850 57052 44850 57052 0 net252
rlabel metal2 46138 56593 46138 56593 0 net253
rlabel metal1 43378 54842 43378 54842 0 net254
rlabel metal1 45172 55930 45172 55930 0 net255
rlabel metal1 46828 57018 46828 57018 0 net256
rlabel metal1 47472 56338 47472 56338 0 net257
rlabel metal1 48852 57018 48852 57018 0 net258
rlabel metal2 23230 56508 23230 56508 0 net26
rlabel metal2 23782 56372 23782 56372 0 net27
rlabel metal2 25898 56304 25898 56304 0 net28
rlabel metal1 30406 57392 30406 57392 0 net29
rlabel metal1 33028 54162 33028 54162 0 net3
rlabel metal1 29302 56678 29302 56678 0 net30
rlabel metal1 10856 57426 10856 57426 0 net31
rlabel metal2 11914 57375 11914 57375 0 net32
rlabel metal2 13294 57596 13294 57596 0 net33
rlabel metal1 14674 57358 14674 57358 0 net34
rlabel via1 21482 57477 21482 57477 0 net35
rlabel metal2 17434 56644 17434 56644 0 net36
rlabel metal1 50278 57018 50278 57018 0 net37
rlabel metal1 51612 57018 51612 57018 0 net38
rlabel metal1 53038 57018 53038 57018 0 net39
rlabel metal2 32430 56542 32430 56542 0 net4
rlabel metal1 54372 57018 54372 57018 0 net40
rlabel metal1 56166 57426 56166 57426 0 net41
rlabel metal1 6532 57018 6532 57018 0 net42
rlabel metal2 8326 57647 8326 57647 0 net43
rlabel metal1 9200 57426 9200 57426 0 net44
rlabel metal1 29900 54842 29900 54842 0 net45
rlabel metal1 31372 54842 31372 54842 0 net46
rlabel metal1 33396 55182 33396 55182 0 net47
rlabel metal1 36110 55114 36110 55114 0 net48
rlabel metal1 37352 55114 37352 55114 0 net49
rlabel metal2 28014 55964 28014 55964 0 net5
rlabel metal2 37306 54706 37306 54706 0 net50
rlabel metal1 38410 54162 38410 54162 0 net51
rlabel metal1 39560 54162 39560 54162 0 net52
rlabel metal2 41078 56372 41078 56372 0 net53
rlabel metal2 46966 56661 46966 56661 0 net54
rlabel metal1 45632 56202 45632 56202 0 net55
rlabel metal1 46000 56338 46000 56338 0 net56
rlabel metal1 47610 56950 47610 56950 0 net57
rlabel metal1 48116 56338 48116 56338 0 net58
rlabel metal2 49726 57120 49726 57120 0 net59
rlabel metal1 34822 55080 34822 55080 0 net6
rlabel metal1 50830 57018 50830 57018 0 net60
rlabel metal2 52486 57222 52486 57222 0 net61
rlabel metal1 53590 57018 53590 57018 0 net62
rlabel metal2 54786 58048 54786 58048 0 net63
rlabel metal1 56212 57018 56212 57018 0 net64
rlabel metal2 17342 1792 17342 1792 0 net65
rlabel metal2 17618 1656 17618 1656 0 net66
rlabel metal2 17894 2132 17894 2132 0 net67
rlabel metal2 18170 1690 18170 1690 0 net68
rlabel metal2 18446 2336 18446 2336 0 net69
rlabel metal1 35604 57426 35604 57426 0 net7
rlabel metal2 18722 2132 18722 2132 0 net70
rlabel metal2 18998 1860 18998 1860 0 net71
rlabel metal2 19274 2132 19274 2132 0 net72
rlabel metal2 19550 1027 19550 1027 0 net73
rlabel metal2 19826 1095 19826 1095 0 net74
rlabel metal2 20102 2336 20102 2336 0 net75
rlabel metal2 20378 2336 20378 2336 0 net76
rlabel metal2 20654 1775 20654 1775 0 net77
rlabel metal2 20930 1792 20930 1792 0 net78
rlabel metal2 21206 2166 21206 2166 0 net79
rlabel metal1 34730 55318 34730 55318 0 net8
rlabel metal2 21482 1554 21482 1554 0 net80
rlabel metal2 21758 2200 21758 2200 0 net81
rlabel metal2 22034 2676 22034 2676 0 net82
rlabel metal1 21666 4046 21666 4046 0 net83
rlabel metal1 22632 4998 22632 4998 0 net84
rlabel metal2 22862 1761 22862 1761 0 net85
rlabel metal2 23138 1656 23138 1656 0 net86
rlabel metal1 23460 5678 23460 5678 0 net87
rlabel metal2 23690 1418 23690 1418 0 net88
rlabel metal1 23184 4726 23184 4726 0 net89
rlabel metal2 34638 57052 34638 57052 0 net9
rlabel metal1 20930 3468 20930 3468 0 net90
rlabel metal1 20194 3026 20194 3026 0 net91
rlabel metal2 24794 1554 24794 1554 0 net92
rlabel metal1 23046 2958 23046 2958 0 net93
rlabel metal2 25346 1384 25346 1384 0 net94
rlabel metal2 25622 1078 25622 1078 0 net95
rlabel metal2 25898 1520 25898 1520 0 net96
rlabel metal2 35006 1367 35006 1367 0 net97
rlabel metal2 35282 959 35282 959 0 net98
rlabel metal1 37812 3366 37812 3366 0 net99
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
