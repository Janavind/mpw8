// This is the unpowered netlist.
module macro_10 (io_active,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input io_active;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net228;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net229;
 wire net257;
 wire net258;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net46;
 wire net47;
 wire net43;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net44;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net45;
 wire net66;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net76;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net77;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net67;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net68;
 wire net96;
 wire net97;
 wire net69;
 wire net70;
 wire net71;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net72;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net73;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net74;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net75;
 wire net162;
 wire net163;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net164;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net165;
 wire net193;
 wire net194;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;

 sky130_fd_sc_hd__clkinv_2 _157_ (.A(net1),
    .Y(_124_));
 sky130_fd_sc_hd__buf_4 _158_ (.A(net1),
    .X(_089_));
 sky130_fd_sc_hd__buf_4 _159_ (.A(_089_),
    .X(_090_));
 sky130_fd_sc_hd__inv_2 _160_ (.A(_090_),
    .Y(_123_));
 sky130_fd_sc_hd__inv_2 _161_ (.A(_090_),
    .Y(_122_));
 sky130_fd_sc_hd__inv_2 _162_ (.A(_090_),
    .Y(_121_));
 sky130_fd_sc_hd__inv_2 _163_ (.A(_090_),
    .Y(_120_));
 sky130_fd_sc_hd__inv_2 _164_ (.A(_090_),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _165_ (.A(_090_),
    .Y(_118_));
 sky130_fd_sc_hd__inv_2 _166_ (.A(_090_),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _167_ (.A(_090_),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _168_ (.A(_090_),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _169_ (.A(_090_),
    .Y(_114_));
 sky130_fd_sc_hd__buf_4 _170_ (.A(_089_),
    .X(_091_));
 sky130_fd_sc_hd__inv_2 _171_ (.A(_091_),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _172_ (.A(_091_),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _173_ (.A(_091_),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _174_ (.A(_091_),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _175_ (.A(_091_),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _176_ (.A(_091_),
    .Y(_108_));
 sky130_fd_sc_hd__inv_2 _177_ (.A(_091_),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _178_ (.A(_091_),
    .Y(_106_));
 sky130_fd_sc_hd__inv_2 _179_ (.A(_091_),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _180_ (.A(_091_),
    .Y(_104_));
 sky130_fd_sc_hd__buf_4 _181_ (.A(_089_),
    .X(_092_));
 sky130_fd_sc_hd__inv_2 _182_ (.A(_092_),
    .Y(_103_));
 sky130_fd_sc_hd__inv_2 _183_ (.A(_092_),
    .Y(_102_));
 sky130_fd_sc_hd__inv_2 _184_ (.A(_092_),
    .Y(_101_));
 sky130_fd_sc_hd__inv_2 _185_ (.A(_092_),
    .Y(_100_));
 sky130_fd_sc_hd__inv_2 _186_ (.A(_092_),
    .Y(_099_));
 sky130_fd_sc_hd__inv_2 _187_ (.A(_092_),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _188_ (.A(_092_),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _189_ (.A(_092_),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _190_ (.A(_092_),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _191_ (.A(_092_),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _192_ (.A(_089_),
    .Y(_093_));
 sky130_fd_sc_hd__nand2b_1 _193_ (.A_N(net19),
    .B(net18),
    .Y(_000_));
 sky130_fd_sc_hd__o31a_1 _194_ (.A1(net8),
    .A2(net6),
    .A3(net7),
    .B1(_000_),
    .X(_001_));
 sky130_fd_sc_hd__xnor2_1 _195_ (.A(net9),
    .B(_001_),
    .Y(_002_));
 sky130_fd_sc_hd__or2_1 _196_ (.A(net5),
    .B(_002_),
    .X(_003_));
 sky130_fd_sc_hd__o21a_1 _197_ (.A1(net6),
    .A2(net7),
    .B1(_000_),
    .X(_004_));
 sky130_fd_sc_hd__xnor2_1 _198_ (.A(net8),
    .B(_004_),
    .Y(_005_));
 sky130_fd_sc_hd__or2_1 _199_ (.A(net4),
    .B(_005_),
    .X(_006_));
 sky130_fd_sc_hd__nand3b_1 _200_ (.A_N(net7),
    .B(_000_),
    .C(net6),
    .Y(_007_));
 sky130_fd_sc_hd__a21bo_1 _201_ (.A1(net6),
    .A2(_000_),
    .B1_N(net7),
    .X(_008_));
 sky130_fd_sc_hd__a21o_1 _202_ (.A1(_007_),
    .A2(_008_),
    .B1(net3),
    .X(_009_));
 sky130_fd_sc_hd__or2b_1 _203_ (.A(net2),
    .B_N(net6),
    .X(_010_));
 sky130_fd_sc_hd__and3_1 _204_ (.A(net3),
    .B(_007_),
    .C(_008_),
    .X(_011_));
 sky130_fd_sc_hd__a21o_1 _205_ (.A1(_009_),
    .A2(_010_),
    .B1(_011_),
    .X(_012_));
 sky130_fd_sc_hd__and2_1 _206_ (.A(net5),
    .B(_002_),
    .X(_013_));
 sky130_fd_sc_hd__and2_1 _207_ (.A(net4),
    .B(_005_),
    .X(_014_));
 sky130_fd_sc_hd__a211o_1 _208_ (.A1(_006_),
    .A2(_012_),
    .B1(_013_),
    .C1(_014_),
    .X(_015_));
 sky130_fd_sc_hd__a21oi_1 _209_ (.A1(net9),
    .A2(_000_),
    .B1(_001_),
    .Y(_016_));
 sky130_fd_sc_hd__a21oi_1 _210_ (.A1(_003_),
    .A2(_015_),
    .B1(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__a31o_1 _211_ (.A1(_016_),
    .A2(_003_),
    .A3(_015_),
    .B1(net19),
    .X(_018_));
 sky130_fd_sc_hd__or2_1 _212_ (.A(_017_),
    .B(_018_),
    .X(_019_));
 sky130_fd_sc_hd__nand2b_1 _213_ (.A_N(net21),
    .B(net20),
    .Y(_020_));
 sky130_fd_sc_hd__o31a_1 _214_ (.A1(net16),
    .A2(net14),
    .A3(net15),
    .B1(_020_),
    .X(_021_));
 sky130_fd_sc_hd__xnor2_1 _215_ (.A(net17),
    .B(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__or2_1 _216_ (.A(net13),
    .B(_022_),
    .X(_023_));
 sky130_fd_sc_hd__o21a_1 _217_ (.A1(net14),
    .A2(net15),
    .B1(_020_),
    .X(_024_));
 sky130_fd_sc_hd__xnor2_1 _218_ (.A(net16),
    .B(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__or2_1 _219_ (.A(net12),
    .B(_025_),
    .X(_026_));
 sky130_fd_sc_hd__nand3b_1 _220_ (.A_N(net15),
    .B(_020_),
    .C(net14),
    .Y(_027_));
 sky130_fd_sc_hd__a21bo_1 _221_ (.A1(net14),
    .A2(_020_),
    .B1_N(net15),
    .X(_028_));
 sky130_fd_sc_hd__a21o_1 _222_ (.A1(_027_),
    .A2(_028_),
    .B1(net11),
    .X(_029_));
 sky130_fd_sc_hd__or2b_1 _223_ (.A(net10),
    .B_N(net14),
    .X(_030_));
 sky130_fd_sc_hd__and3_1 _224_ (.A(net11),
    .B(_027_),
    .C(_028_),
    .X(_031_));
 sky130_fd_sc_hd__a21o_1 _225_ (.A1(_029_),
    .A2(_030_),
    .B1(_031_),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _226_ (.A(net13),
    .B(_022_),
    .X(_033_));
 sky130_fd_sc_hd__and2_1 _227_ (.A(net12),
    .B(_025_),
    .X(_034_));
 sky130_fd_sc_hd__a211o_1 _228_ (.A1(_026_),
    .A2(_032_),
    .B1(_033_),
    .C1(_034_),
    .X(_035_));
 sky130_fd_sc_hd__a21oi_1 _229_ (.A1(net17),
    .A2(_020_),
    .B1(_021_),
    .Y(_036_));
 sky130_fd_sc_hd__a21oi_1 _230_ (.A1(_023_),
    .A2(_035_),
    .B1(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__a31o_1 _231_ (.A1(_036_),
    .A2(_023_),
    .A3(_035_),
    .B1(net21),
    .X(_038_));
 sky130_fd_sc_hd__or2_1 _232_ (.A(_037_),
    .B(_038_),
    .X(_039_));
 sky130_fd_sc_hd__nor3_2 _233_ (.A(_124_),
    .B(_037_),
    .C(_038_),
    .Y(net31));
 sky130_fd_sc_hd__nor3_1 _234_ (.A(_124_),
    .B(_017_),
    .C(_018_),
    .Y(net32));
 sky130_fd_sc_hd__o22a_1 _235_ (.A1(_019_),
    .A2(_039_),
    .B1(net31),
    .B2(net32),
    .X(net22));
 sky130_fd_sc_hd__inv_2 _236_ (.A(net19),
    .Y(_040_));
 sky130_fd_sc_hd__o2bb2a_1 _237_ (.A1_N(net6),
    .A2_N(net2),
    .B1(_040_),
    .B2(net18),
    .X(_041_));
 sky130_fd_sc_hd__o21a_1 _238_ (.A1(net6),
    .A2(net2),
    .B1(_041_),
    .X(_042_));
 sky130_fd_sc_hd__a31o_1 _239_ (.A1(net6),
    .A2(net19),
    .A3(net2),
    .B1(_042_),
    .X(_043_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(net21),
    .Y(_044_));
 sky130_fd_sc_hd__o2bb2a_1 _241_ (.A1_N(net14),
    .A2_N(net10),
    .B1(_044_),
    .B2(net20),
    .X(_045_));
 sky130_fd_sc_hd__o21a_1 _242_ (.A1(net14),
    .A2(net10),
    .B1(_045_),
    .X(_046_));
 sky130_fd_sc_hd__a31o_1 _243_ (.A1(net14),
    .A2(net21),
    .A3(net10),
    .B1(_046_),
    .X(_047_));
 sky130_fd_sc_hd__and2_1 _244_ (.A(_089_),
    .B(_047_),
    .X(_048_));
 sky130_fd_sc_hd__clkbuf_1 _245_ (.A(_048_),
    .X(net23));
 sky130_fd_sc_hd__and2_1 _246_ (.A(_089_),
    .B(_043_),
    .X(_049_));
 sky130_fd_sc_hd__clkbuf_1 _247_ (.A(_049_),
    .X(net27));
 sky130_fd_sc_hd__o2bb2a_1 _248_ (.A1_N(_043_),
    .A2_N(_047_),
    .B1(net23),
    .B2(net27),
    .X(net33));
 sky130_fd_sc_hd__or2b_1 _249_ (.A(_011_),
    .B_N(_009_),
    .X(_050_));
 sky130_fd_sc_hd__xnor2_1 _250_ (.A(_050_),
    .B(_010_),
    .Y(_051_));
 sky130_fd_sc_hd__o21a_1 _251_ (.A1(net7),
    .A2(net18),
    .B1(net3),
    .X(_052_));
 sky130_fd_sc_hd__a211o_1 _252_ (.A1(net7),
    .A2(net18),
    .B1(_040_),
    .C1(_052_),
    .X(_053_));
 sky130_fd_sc_hd__o21a_1 _253_ (.A1(net19),
    .A2(_051_),
    .B1(_053_),
    .X(_054_));
 sky130_fd_sc_hd__or2b_1 _254_ (.A(_031_),
    .B_N(_029_),
    .X(_055_));
 sky130_fd_sc_hd__xnor2_1 _255_ (.A(_055_),
    .B(_030_),
    .Y(_056_));
 sky130_fd_sc_hd__o21a_1 _256_ (.A1(net15),
    .A2(net20),
    .B1(net11),
    .X(_057_));
 sky130_fd_sc_hd__a211o_1 _257_ (.A1(net15),
    .A2(net20),
    .B1(_044_),
    .C1(_057_),
    .X(_058_));
 sky130_fd_sc_hd__o21a_1 _258_ (.A1(net21),
    .A2(_056_),
    .B1(_058_),
    .X(_059_));
 sky130_fd_sc_hd__and2_1 _259_ (.A(_089_),
    .B(_059_),
    .X(_060_));
 sky130_fd_sc_hd__clkbuf_1 _260_ (.A(_060_),
    .X(net24));
 sky130_fd_sc_hd__and2_1 _261_ (.A(_089_),
    .B(_054_),
    .X(_061_));
 sky130_fd_sc_hd__clkbuf_1 _262_ (.A(_061_),
    .X(net28));
 sky130_fd_sc_hd__o2bb2a_1 _263_ (.A1_N(_054_),
    .A2_N(_059_),
    .B1(net24),
    .B2(net28),
    .X(net34));
 sky130_fd_sc_hd__a21o_1 _264_ (.A1(net18),
    .A2(net4),
    .B1(net8),
    .X(_062_));
 sky130_fd_sc_hd__or2_1 _265_ (.A(net18),
    .B(net4),
    .X(_063_));
 sky130_fd_sc_hd__xor2_1 _266_ (.A(net4),
    .B(_005_),
    .X(_064_));
 sky130_fd_sc_hd__or2_1 _267_ (.A(_064_),
    .B(_012_),
    .X(_065_));
 sky130_fd_sc_hd__a21oi_1 _268_ (.A1(_064_),
    .A2(_012_),
    .B1(net19),
    .Y(_066_));
 sky130_fd_sc_hd__a32o_1 _269_ (.A1(net19),
    .A2(_062_),
    .A3(_063_),
    .B1(_065_),
    .B2(_066_),
    .X(_067_));
 sky130_fd_sc_hd__a21o_1 _270_ (.A1(net20),
    .A2(net12),
    .B1(net16),
    .X(_068_));
 sky130_fd_sc_hd__or2_1 _271_ (.A(net20),
    .B(net12),
    .X(_069_));
 sky130_fd_sc_hd__xor2_1 _272_ (.A(net12),
    .B(_025_),
    .X(_070_));
 sky130_fd_sc_hd__or2_1 _273_ (.A(_070_),
    .B(_032_),
    .X(_071_));
 sky130_fd_sc_hd__a21oi_1 _274_ (.A1(_070_),
    .A2(_032_),
    .B1(net21),
    .Y(_072_));
 sky130_fd_sc_hd__a32o_1 _275_ (.A1(net21),
    .A2(_068_),
    .A3(_069_),
    .B1(_071_),
    .B2(_072_),
    .X(_073_));
 sky130_fd_sc_hd__and2_1 _276_ (.A(net1),
    .B(_073_),
    .X(_074_));
 sky130_fd_sc_hd__clkbuf_1 _277_ (.A(_074_),
    .X(net25));
 sky130_fd_sc_hd__and2_1 _278_ (.A(_089_),
    .B(_067_),
    .X(_075_));
 sky130_fd_sc_hd__clkbuf_1 _279_ (.A(_075_),
    .X(net29));
 sky130_fd_sc_hd__o2bb2a_1 _280_ (.A1_N(_067_),
    .A2_N(_073_),
    .B1(net25),
    .B2(net29),
    .X(net35));
 sky130_fd_sc_hd__a21oi_1 _281_ (.A1(_006_),
    .A2(_012_),
    .B1(_014_),
    .Y(_076_));
 sky130_fd_sc_hd__and2b_1 _282_ (.A_N(_013_),
    .B(_003_),
    .X(_077_));
 sky130_fd_sc_hd__xnor2_1 _283_ (.A(_076_),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__nor2_1 _284_ (.A(net19),
    .B(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__o21a_1 _285_ (.A1(net9),
    .A2(net18),
    .B1(net5),
    .X(_080_));
 sky130_fd_sc_hd__a21o_1 _286_ (.A1(net9),
    .A2(net18),
    .B1(_040_),
    .X(_081_));
 sky130_fd_sc_hd__nor2_1 _287_ (.A(_080_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__a21o_1 _288_ (.A1(_026_),
    .A2(_032_),
    .B1(_034_),
    .X(_083_));
 sky130_fd_sc_hd__and2b_1 _289_ (.A_N(_033_),
    .B(_023_),
    .X(_084_));
 sky130_fd_sc_hd__xnor2_1 _290_ (.A(_083_),
    .B(_084_),
    .Y(_085_));
 sky130_fd_sc_hd__o21a_1 _291_ (.A1(net17),
    .A2(net20),
    .B1(net13),
    .X(_086_));
 sky130_fd_sc_hd__a211oi_2 _292_ (.A1(net17),
    .A2(net20),
    .B1(_044_),
    .C1(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__a21o_1 _293_ (.A1(_044_),
    .A2(_085_),
    .B1(_087_),
    .X(_088_));
 sky130_fd_sc_hd__a211oi_2 _294_ (.A1(_044_),
    .A2(_085_),
    .B1(_087_),
    .C1(_124_),
    .Y(net26));
 sky130_fd_sc_hd__o221a_1 _295_ (.A1(net19),
    .A2(_078_),
    .B1(_080_),
    .B2(_081_),
    .C1(_089_),
    .X(net30));
 sky130_fd_sc_hd__o32a_1 _296_ (.A1(_079_),
    .A2(_082_),
    .A3(_088_),
    .B1(net26),
    .B2(net30),
    .X(net36));
 sky130_fd_sc_hd__conb_1 macro_10_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 macro_10_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 macro_10_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 macro_10_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 macro_10_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 macro_10_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 macro_10_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 macro_10_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 macro_10_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 macro_10_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 macro_10_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 macro_10_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 macro_10_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 macro_10_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 macro_10_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 macro_10_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 macro_10_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 macro_10_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 macro_10_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 macro_10_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 macro_10_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 macro_10_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 macro_10_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 macro_10_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 macro_10_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 macro_10_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 macro_10_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 macro_10_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 macro_10_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 macro_10_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 macro_10_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 macro_10_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 macro_10_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 macro_10_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 macro_10_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 macro_10_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 macro_10_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 macro_10_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 macro_10_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 macro_10_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 macro_10_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 macro_10_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 macro_10_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 macro_10_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 macro_10_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 macro_10_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 macro_10_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 macro_10_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 macro_10_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 macro_10_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 macro_10_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 macro_10_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 macro_10_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 macro_10_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 macro_10_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 macro_10_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 macro_10_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 macro_10_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 macro_10_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 macro_10_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 macro_10_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 macro_10_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 macro_10_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 macro_10_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 macro_10_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 macro_10_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 macro_10_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 macro_10_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 macro_10_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 macro_10_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 macro_10_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 macro_10_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 macro_10_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 macro_10_111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 macro_10_112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 macro_10_113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 macro_10_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 macro_10_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 macro_10_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 macro_10_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 macro_10_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 macro_10_119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 macro_10_120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 macro_10_121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 macro_10_122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 macro_10_123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 macro_10_124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 macro_10_125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 macro_10_126 (.LO(net126));
 sky130_fd_sc_hd__conb_1 macro_10_127 (.LO(net127));
 sky130_fd_sc_hd__conb_1 macro_10_128 (.LO(net128));
 sky130_fd_sc_hd__conb_1 macro_10_129 (.LO(net129));
 sky130_fd_sc_hd__conb_1 macro_10_130 (.LO(net130));
 sky130_fd_sc_hd__conb_1 macro_10_131 (.LO(net131));
 sky130_fd_sc_hd__conb_1 macro_10_132 (.LO(net132));
 sky130_fd_sc_hd__conb_1 macro_10_133 (.LO(net133));
 sky130_fd_sc_hd__conb_1 macro_10_134 (.LO(net134));
 sky130_fd_sc_hd__conb_1 macro_10_135 (.LO(net135));
 sky130_fd_sc_hd__conb_1 macro_10_136 (.LO(net136));
 sky130_fd_sc_hd__conb_1 macro_10_137 (.LO(net137));
 sky130_fd_sc_hd__conb_1 macro_10_138 (.LO(net138));
 sky130_fd_sc_hd__conb_1 macro_10_139 (.LO(net139));
 sky130_fd_sc_hd__conb_1 macro_10_140 (.LO(net140));
 sky130_fd_sc_hd__conb_1 macro_10_141 (.LO(net141));
 sky130_fd_sc_hd__conb_1 macro_10_142 (.LO(net142));
 sky130_fd_sc_hd__conb_1 macro_10_143 (.LO(net143));
 sky130_fd_sc_hd__conb_1 macro_10_144 (.LO(net144));
 sky130_fd_sc_hd__conb_1 macro_10_145 (.LO(net145));
 sky130_fd_sc_hd__conb_1 macro_10_146 (.LO(net146));
 sky130_fd_sc_hd__conb_1 macro_10_147 (.LO(net147));
 sky130_fd_sc_hd__conb_1 macro_10_148 (.LO(net148));
 sky130_fd_sc_hd__conb_1 macro_10_149 (.LO(net149));
 sky130_fd_sc_hd__conb_1 macro_10_150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 macro_10_151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 macro_10_152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 macro_10_153 (.LO(net153));
 sky130_fd_sc_hd__conb_1 macro_10_154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 macro_10_155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 macro_10_156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 macro_10_157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 macro_10_158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 macro_10_159 (.LO(net159));
 sky130_fd_sc_hd__conb_1 macro_10_160 (.LO(net160));
 sky130_fd_sc_hd__conb_1 macro_10_161 (.LO(net161));
 sky130_fd_sc_hd__conb_1 macro_10_162 (.LO(net162));
 sky130_fd_sc_hd__conb_1 macro_10_163 (.LO(net163));
 sky130_fd_sc_hd__conb_1 macro_10_164 (.LO(net164));
 sky130_fd_sc_hd__conb_1 macro_10_165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 macro_10_166 (.LO(net166));
 sky130_fd_sc_hd__conb_1 macro_10_167 (.LO(net167));
 sky130_fd_sc_hd__conb_1 macro_10_168 (.LO(net168));
 sky130_fd_sc_hd__conb_1 macro_10_169 (.LO(net169));
 sky130_fd_sc_hd__conb_1 macro_10_170 (.LO(net170));
 sky130_fd_sc_hd__conb_1 macro_10_171 (.LO(net171));
 sky130_fd_sc_hd__conb_1 macro_10_172 (.LO(net172));
 sky130_fd_sc_hd__conb_1 macro_10_173 (.LO(net173));
 sky130_fd_sc_hd__conb_1 macro_10_174 (.LO(net174));
 sky130_fd_sc_hd__conb_1 macro_10_175 (.LO(net175));
 sky130_fd_sc_hd__conb_1 macro_10_176 (.LO(net176));
 sky130_fd_sc_hd__conb_1 macro_10_177 (.LO(net177));
 sky130_fd_sc_hd__conb_1 macro_10_178 (.LO(net178));
 sky130_fd_sc_hd__conb_1 macro_10_179 (.LO(net179));
 sky130_fd_sc_hd__conb_1 macro_10_180 (.LO(net180));
 sky130_fd_sc_hd__conb_1 macro_10_181 (.LO(net181));
 sky130_fd_sc_hd__conb_1 macro_10_182 (.LO(net182));
 sky130_fd_sc_hd__conb_1 macro_10_183 (.LO(net183));
 sky130_fd_sc_hd__conb_1 macro_10_184 (.LO(net184));
 sky130_fd_sc_hd__conb_1 macro_10_185 (.LO(net185));
 sky130_fd_sc_hd__conb_1 macro_10_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 macro_10_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 macro_10_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 macro_10_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 macro_10_190 (.LO(net190));
 sky130_fd_sc_hd__conb_1 macro_10_191 (.LO(net191));
 sky130_fd_sc_hd__conb_1 macro_10_192 (.LO(net192));
 sky130_fd_sc_hd__conb_1 macro_10_193 (.LO(net193));
 sky130_fd_sc_hd__conb_1 _519__194 (.LO(net194));
 sky130_fd_sc_hd__conb_1 _520__195 (.LO(net195));
 sky130_fd_sc_hd__conb_1 _521__196 (.LO(net196));
 sky130_fd_sc_hd__conb_1 _522__197 (.LO(net197));
 sky130_fd_sc_hd__conb_1 _523__198 (.LO(net198));
 sky130_fd_sc_hd__conb_1 _524__199 (.LO(net199));
 sky130_fd_sc_hd__conb_1 _525__200 (.LO(net200));
 sky130_fd_sc_hd__conb_1 _526__201 (.LO(net201));
 sky130_fd_sc_hd__conb_1 _527__202 (.LO(net202));
 sky130_fd_sc_hd__conb_1 _528__203 (.LO(net203));
 sky130_fd_sc_hd__conb_1 _529__204 (.LO(net204));
 sky130_fd_sc_hd__conb_1 _530__205 (.LO(net205));
 sky130_fd_sc_hd__conb_1 _531__206 (.LO(net206));
 sky130_fd_sc_hd__conb_1 _532__207 (.LO(net207));
 sky130_fd_sc_hd__conb_1 _533__208 (.LO(net208));
 sky130_fd_sc_hd__conb_1 _534__209 (.LO(net209));
 sky130_fd_sc_hd__conb_1 _535__210 (.LO(net210));
 sky130_fd_sc_hd__conb_1 _536__211 (.LO(net211));
 sky130_fd_sc_hd__conb_1 _537__212 (.LO(net212));
 sky130_fd_sc_hd__conb_1 _538__213 (.LO(net213));
 sky130_fd_sc_hd__conb_1 _539__214 (.LO(net214));
 sky130_fd_sc_hd__conb_1 _540__215 (.LO(net215));
 sky130_fd_sc_hd__conb_1 _541__216 (.LO(net216));
 sky130_fd_sc_hd__conb_1 _542__217 (.LO(net217));
 sky130_fd_sc_hd__conb_1 _543__218 (.LO(net218));
 sky130_fd_sc_hd__conb_1 _544__219 (.LO(net219));
 sky130_fd_sc_hd__conb_1 _545__220 (.LO(net220));
 sky130_fd_sc_hd__conb_1 _546__221 (.LO(net221));
 sky130_fd_sc_hd__conb_1 _547__222 (.LO(net222));
 sky130_fd_sc_hd__conb_1 _548__223 (.LO(net223));
 sky130_fd_sc_hd__conb_1 _549__224 (.LO(net224));
 sky130_fd_sc_hd__conb_1 _550__225 (.LO(net225));
 sky130_fd_sc_hd__conb_1 macro_10_226 (.LO(net226));
 sky130_fd_sc_hd__conb_1 macro_10_227 (.LO(net227));
 sky130_fd_sc_hd__conb_1 macro_10_228 (.LO(net228));
 sky130_fd_sc_hd__conb_1 macro_10_229 (.LO(net229));
 sky130_fd_sc_hd__conb_1 macro_10_230 (.LO(net230));
 sky130_fd_sc_hd__conb_1 macro_10_231 (.LO(net231));
 sky130_fd_sc_hd__conb_1 macro_10_232 (.LO(net232));
 sky130_fd_sc_hd__conb_1 macro_10_233 (.LO(net233));
 sky130_fd_sc_hd__conb_1 macro_10_234 (.LO(net234));
 sky130_fd_sc_hd__conb_1 macro_10_235 (.LO(net235));
 sky130_fd_sc_hd__conb_1 macro_10_236 (.LO(net236));
 sky130_fd_sc_hd__conb_1 macro_10_237 (.LO(net237));
 sky130_fd_sc_hd__conb_1 macro_10_238 (.LO(net238));
 sky130_fd_sc_hd__conb_1 macro_10_239 (.LO(net239));
 sky130_fd_sc_hd__conb_1 macro_10_240 (.LO(net240));
 sky130_fd_sc_hd__conb_1 macro_10_241 (.LO(net241));
 sky130_fd_sc_hd__conb_1 macro_10_242 (.LO(net242));
 sky130_fd_sc_hd__conb_1 macro_10_243 (.LO(net243));
 sky130_fd_sc_hd__conb_1 macro_10_244 (.LO(net244));
 sky130_fd_sc_hd__conb_1 macro_10_245 (.LO(net245));
 sky130_fd_sc_hd__conb_1 macro_10_246 (.LO(net246));
 sky130_fd_sc_hd__conb_1 macro_10_247 (.LO(net247));
 sky130_fd_sc_hd__conb_1 macro_10_248 (.LO(net248));
 sky130_fd_sc_hd__conb_1 macro_10_249 (.LO(net249));
 sky130_fd_sc_hd__conb_1 macro_10_250 (.LO(net250));
 sky130_fd_sc_hd__conb_1 macro_10_251 (.LO(net251));
 sky130_fd_sc_hd__conb_1 macro_10_252 (.LO(net252));
 sky130_fd_sc_hd__conb_1 macro_10_253 (.LO(net253));
 sky130_fd_sc_hd__conb_1 macro_10_254 (.LO(net254));
 sky130_fd_sc_hd__conb_1 macro_10_255 (.LO(net255));
 sky130_fd_sc_hd__conb_1 macro_10_256 (.LO(net256));
 sky130_fd_sc_hd__conb_1 macro_10_257 (.LO(net257));
 sky130_fd_sc_hd__conb_1 macro_10_258 (.LO(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__C1 (.DIODE(_089_));
 sky130_fd_sc_hd__ebufn_8 _519_ (.A(net194),
    .TE_B(_093_),
    .Z(la_data_out[32]));
 sky130_fd_sc_hd__ebufn_8 _520_ (.A(net195),
    .TE_B(_094_),
    .Z(la_data_out[33]));
 sky130_fd_sc_hd__ebufn_8 _521_ (.A(net196),
    .TE_B(_095_),
    .Z(la_data_out[34]));
 sky130_fd_sc_hd__ebufn_8 _522_ (.A(net197),
    .TE_B(_096_),
    .Z(la_data_out[35]));
 sky130_fd_sc_hd__ebufn_8 _523_ (.A(net198),
    .TE_B(_097_),
    .Z(la_data_out[36]));
 sky130_fd_sc_hd__ebufn_8 _524_ (.A(net199),
    .TE_B(_098_),
    .Z(la_data_out[37]));
 sky130_fd_sc_hd__ebufn_8 _525_ (.A(net200),
    .TE_B(_099_),
    .Z(la_data_out[38]));
 sky130_fd_sc_hd__ebufn_8 _526_ (.A(net201),
    .TE_B(_100_),
    .Z(la_data_out[39]));
 sky130_fd_sc_hd__ebufn_8 _527_ (.A(net202),
    .TE_B(_101_),
    .Z(la_data_out[40]));
 sky130_fd_sc_hd__ebufn_8 _528_ (.A(net203),
    .TE_B(_102_),
    .Z(la_data_out[41]));
 sky130_fd_sc_hd__ebufn_8 _529_ (.A(net204),
    .TE_B(_103_),
    .Z(la_data_out[42]));
 sky130_fd_sc_hd__ebufn_8 _530_ (.A(net205),
    .TE_B(_104_),
    .Z(la_data_out[43]));
 sky130_fd_sc_hd__ebufn_8 _531_ (.A(net206),
    .TE_B(_105_),
    .Z(la_data_out[44]));
 sky130_fd_sc_hd__ebufn_8 _532_ (.A(net207),
    .TE_B(_106_),
    .Z(la_data_out[45]));
 sky130_fd_sc_hd__ebufn_8 _533_ (.A(net208),
    .TE_B(_107_),
    .Z(la_data_out[46]));
 sky130_fd_sc_hd__ebufn_8 _534_ (.A(net209),
    .TE_B(_108_),
    .Z(la_data_out[47]));
 sky130_fd_sc_hd__ebufn_8 _535_ (.A(net210),
    .TE_B(_109_),
    .Z(la_data_out[48]));
 sky130_fd_sc_hd__ebufn_8 _536_ (.A(net211),
    .TE_B(_110_),
    .Z(la_data_out[49]));
 sky130_fd_sc_hd__ebufn_8 _537_ (.A(net212),
    .TE_B(_111_),
    .Z(la_data_out[50]));
 sky130_fd_sc_hd__ebufn_8 _538_ (.A(net213),
    .TE_B(_112_),
    .Z(la_data_out[51]));
 sky130_fd_sc_hd__ebufn_8 _539_ (.A(net214),
    .TE_B(_113_),
    .Z(la_data_out[52]));
 sky130_fd_sc_hd__ebufn_8 _540_ (.A(net215),
    .TE_B(_114_),
    .Z(la_data_out[53]));
 sky130_fd_sc_hd__ebufn_8 _541_ (.A(net216),
    .TE_B(_115_),
    .Z(la_data_out[54]));
 sky130_fd_sc_hd__ebufn_8 _542_ (.A(net217),
    .TE_B(_116_),
    .Z(la_data_out[55]));
 sky130_fd_sc_hd__ebufn_8 _543_ (.A(net218),
    .TE_B(_117_),
    .Z(la_data_out[56]));
 sky130_fd_sc_hd__ebufn_8 _544_ (.A(net219),
    .TE_B(_118_),
    .Z(la_data_out[57]));
 sky130_fd_sc_hd__ebufn_8 _545_ (.A(net220),
    .TE_B(_119_),
    .Z(la_data_out[58]));
 sky130_fd_sc_hd__ebufn_8 _546_ (.A(net221),
    .TE_B(_120_),
    .Z(la_data_out[59]));
 sky130_fd_sc_hd__ebufn_8 _547_ (.A(net222),
    .TE_B(_121_),
    .Z(la_data_out[60]));
 sky130_fd_sc_hd__ebufn_8 _548_ (.A(net223),
    .TE_B(_122_),
    .Z(la_data_out[61]));
 sky130_fd_sc_hd__ebufn_8 _549_ (.A(net224),
    .TE_B(_123_),
    .Z(la_data_out[62]));
 sky130_fd_sc_hd__ebufn_8 _550_ (.A(net225),
    .TE_B(_124_),
    .Z(la_data_out[63]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_active),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[18]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[19]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(io_in[20]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[21]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[22]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(io_in[23]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(io_in[24]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(io_in[25]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(io_in[26]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(io_in[27]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(io_in[28]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(io_in[29]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(io_in[30]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(io_in[31]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(io_in[32]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(io_in[33]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(io_in[34]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(io_in[35]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(io_in[36]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(io_in[37]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(io_out[9]));
 sky130_fd_sc_hd__conb_1 macro_10_37 (.LO(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__278__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__261__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__259__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__246__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__170__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__159__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_active));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(io_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(io_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(io_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__157__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__286__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__285__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__265__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__284__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__269__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__253__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__236__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__A_N (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__274__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__231__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__A_N (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__B1 (.DIODE(net31));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_622 ();
 assign io_oeb[0] = net226;
 assign io_oeb[10] = net236;
 assign io_oeb[11] = net237;
 assign io_oeb[12] = net238;
 assign io_oeb[13] = net239;
 assign io_oeb[14] = net240;
 assign io_oeb[15] = net241;
 assign io_oeb[16] = net242;
 assign io_oeb[17] = net243;
 assign io_oeb[18] = net244;
 assign io_oeb[19] = net245;
 assign io_oeb[1] = net227;
 assign io_oeb[20] = net246;
 assign io_oeb[21] = net247;
 assign io_oeb[22] = net248;
 assign io_oeb[23] = net249;
 assign io_oeb[24] = net250;
 assign io_oeb[25] = net251;
 assign io_oeb[26] = net252;
 assign io_oeb[27] = net253;
 assign io_oeb[28] = net254;
 assign io_oeb[29] = net255;
 assign io_oeb[2] = net228;
 assign io_oeb[30] = net256;
 assign io_oeb[31] = net257;
 assign io_oeb[32] = net258;
 assign io_oeb[33] = net37;
 assign io_oeb[34] = net38;
 assign io_oeb[35] = net39;
 assign io_oeb[36] = net40;
 assign io_oeb[37] = net41;
 assign io_oeb[3] = net229;
 assign io_oeb[4] = net230;
 assign io_oeb[5] = net231;
 assign io_oeb[6] = net232;
 assign io_oeb[7] = net233;
 assign io_oeb[8] = net234;
 assign io_oeb[9] = net235;
 assign io_out[18] = net45;
 assign io_out[19] = net46;
 assign io_out[1] = net42;
 assign io_out[20] = net47;
 assign io_out[21] = net48;
 assign io_out[22] = net49;
 assign io_out[23] = net50;
 assign io_out[24] = net51;
 assign io_out[25] = net52;
 assign io_out[26] = net53;
 assign io_out[27] = net54;
 assign io_out[28] = net55;
 assign io_out[29] = net56;
 assign io_out[2] = net43;
 assign io_out[30] = net57;
 assign io_out[31] = net58;
 assign io_out[32] = net59;
 assign io_out[33] = net60;
 assign io_out[34] = net61;
 assign io_out[35] = net62;
 assign io_out[36] = net63;
 assign io_out[37] = net64;
 assign io_out[3] = net44;
 assign la_data_out[0] = net65;
 assign la_data_out[100] = net133;
 assign la_data_out[101] = net134;
 assign la_data_out[102] = net135;
 assign la_data_out[103] = net136;
 assign la_data_out[104] = net137;
 assign la_data_out[105] = net138;
 assign la_data_out[106] = net139;
 assign la_data_out[107] = net140;
 assign la_data_out[108] = net141;
 assign la_data_out[109] = net142;
 assign la_data_out[10] = net75;
 assign la_data_out[110] = net143;
 assign la_data_out[111] = net144;
 assign la_data_out[112] = net145;
 assign la_data_out[113] = net146;
 assign la_data_out[114] = net147;
 assign la_data_out[115] = net148;
 assign la_data_out[116] = net149;
 assign la_data_out[117] = net150;
 assign la_data_out[118] = net151;
 assign la_data_out[119] = net152;
 assign la_data_out[11] = net76;
 assign la_data_out[120] = net153;
 assign la_data_out[121] = net154;
 assign la_data_out[122] = net155;
 assign la_data_out[123] = net156;
 assign la_data_out[124] = net157;
 assign la_data_out[125] = net158;
 assign la_data_out[126] = net159;
 assign la_data_out[127] = net160;
 assign la_data_out[12] = net77;
 assign la_data_out[13] = net78;
 assign la_data_out[14] = net79;
 assign la_data_out[15] = net80;
 assign la_data_out[16] = net81;
 assign la_data_out[17] = net82;
 assign la_data_out[18] = net83;
 assign la_data_out[19] = net84;
 assign la_data_out[1] = net66;
 assign la_data_out[20] = net85;
 assign la_data_out[21] = net86;
 assign la_data_out[22] = net87;
 assign la_data_out[23] = net88;
 assign la_data_out[24] = net89;
 assign la_data_out[25] = net90;
 assign la_data_out[26] = net91;
 assign la_data_out[27] = net92;
 assign la_data_out[28] = net93;
 assign la_data_out[29] = net94;
 assign la_data_out[2] = net67;
 assign la_data_out[30] = net95;
 assign la_data_out[31] = net96;
 assign la_data_out[3] = net68;
 assign la_data_out[4] = net69;
 assign la_data_out[5] = net70;
 assign la_data_out[64] = net97;
 assign la_data_out[65] = net98;
 assign la_data_out[66] = net99;
 assign la_data_out[67] = net100;
 assign la_data_out[68] = net101;
 assign la_data_out[69] = net102;
 assign la_data_out[6] = net71;
 assign la_data_out[70] = net103;
 assign la_data_out[71] = net104;
 assign la_data_out[72] = net105;
 assign la_data_out[73] = net106;
 assign la_data_out[74] = net107;
 assign la_data_out[75] = net108;
 assign la_data_out[76] = net109;
 assign la_data_out[77] = net110;
 assign la_data_out[78] = net111;
 assign la_data_out[79] = net112;
 assign la_data_out[7] = net72;
 assign la_data_out[80] = net113;
 assign la_data_out[81] = net114;
 assign la_data_out[82] = net115;
 assign la_data_out[83] = net116;
 assign la_data_out[84] = net117;
 assign la_data_out[85] = net118;
 assign la_data_out[86] = net119;
 assign la_data_out[87] = net120;
 assign la_data_out[88] = net121;
 assign la_data_out[89] = net122;
 assign la_data_out[8] = net73;
 assign la_data_out[90] = net123;
 assign la_data_out[91] = net124;
 assign la_data_out[92] = net125;
 assign la_data_out[93] = net126;
 assign la_data_out[94] = net127;
 assign la_data_out[95] = net128;
 assign la_data_out[96] = net129;
 assign la_data_out[97] = net130;
 assign la_data_out[98] = net131;
 assign la_data_out[99] = net132;
 assign la_data_out[9] = net74;
 assign wbs_ack_o = net161;
 assign wbs_dat_o[0] = net162;
 assign wbs_dat_o[10] = net172;
 assign wbs_dat_o[11] = net173;
 assign wbs_dat_o[12] = net174;
 assign wbs_dat_o[13] = net175;
 assign wbs_dat_o[14] = net176;
 assign wbs_dat_o[15] = net177;
 assign wbs_dat_o[16] = net178;
 assign wbs_dat_o[17] = net179;
 assign wbs_dat_o[18] = net180;
 assign wbs_dat_o[19] = net181;
 assign wbs_dat_o[1] = net163;
 assign wbs_dat_o[20] = net182;
 assign wbs_dat_o[21] = net183;
 assign wbs_dat_o[22] = net184;
 assign wbs_dat_o[23] = net185;
 assign wbs_dat_o[24] = net186;
 assign wbs_dat_o[25] = net187;
 assign wbs_dat_o[26] = net188;
 assign wbs_dat_o[27] = net189;
 assign wbs_dat_o[28] = net190;
 assign wbs_dat_o[29] = net191;
 assign wbs_dat_o[2] = net164;
 assign wbs_dat_o[30] = net192;
 assign wbs_dat_o[31] = net193;
 assign wbs_dat_o[3] = net165;
 assign wbs_dat_o[4] = net166;
 assign wbs_dat_o[5] = net167;
 assign wbs_dat_o[6] = net168;
 assign wbs_dat_o[7] = net169;
 assign wbs_dat_o[8] = net170;
 assign wbs_dat_o[9] = net171;
endmodule

