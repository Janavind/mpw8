// This is the unpowered netlist.
module macro_decap_12 (io_active,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input io_active;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net228;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net229;
 wire net257;
 wire net258;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net46;
 wire net47;
 wire net43;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net44;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net45;
 wire net66;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net76;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net77;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net67;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net68;
 wire net96;
 wire net97;
 wire net69;
 wire net70;
 wire net71;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net72;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net73;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net74;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net75;
 wire net162;
 wire net163;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net164;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net165;
 wire net193;
 wire net194;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;

 sky130_fd_sc_hd__inv_2 _157_ (.A(net1),
    .Y(_124_));
 sky130_fd_sc_hd__buf_4 _158_ (.A(net1),
    .X(_089_));
 sky130_fd_sc_hd__buf_4 _159_ (.A(_089_),
    .X(_090_));
 sky130_fd_sc_hd__inv_2 _160_ (.A(_090_),
    .Y(_123_));
 sky130_fd_sc_hd__inv_2 _161_ (.A(_090_),
    .Y(_122_));
 sky130_fd_sc_hd__inv_2 _162_ (.A(_090_),
    .Y(_121_));
 sky130_fd_sc_hd__inv_2 _163_ (.A(_090_),
    .Y(_120_));
 sky130_fd_sc_hd__inv_2 _164_ (.A(_090_),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _165_ (.A(_090_),
    .Y(_118_));
 sky130_fd_sc_hd__inv_2 _166_ (.A(_090_),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _167_ (.A(_090_),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _168_ (.A(_090_),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _169_ (.A(_090_),
    .Y(_114_));
 sky130_fd_sc_hd__buf_4 _170_ (.A(_089_),
    .X(_091_));
 sky130_fd_sc_hd__inv_2 _171_ (.A(_091_),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _172_ (.A(_091_),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _173_ (.A(_091_),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _174_ (.A(_091_),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _175_ (.A(_091_),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _176_ (.A(_091_),
    .Y(_108_));
 sky130_fd_sc_hd__inv_2 _177_ (.A(_091_),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _178_ (.A(_091_),
    .Y(_106_));
 sky130_fd_sc_hd__inv_2 _179_ (.A(_091_),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _180_ (.A(_091_),
    .Y(_104_));
 sky130_fd_sc_hd__buf_4 _181_ (.A(_089_),
    .X(_092_));
 sky130_fd_sc_hd__inv_2 _182_ (.A(_092_),
    .Y(_103_));
 sky130_fd_sc_hd__inv_2 _183_ (.A(_092_),
    .Y(_102_));
 sky130_fd_sc_hd__inv_2 _184_ (.A(_092_),
    .Y(_101_));
 sky130_fd_sc_hd__inv_2 _185_ (.A(_092_),
    .Y(_100_));
 sky130_fd_sc_hd__inv_2 _186_ (.A(_092_),
    .Y(_099_));
 sky130_fd_sc_hd__inv_2 _187_ (.A(_092_),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _188_ (.A(_092_),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _189_ (.A(_092_),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _190_ (.A(_092_),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _191_ (.A(_092_),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _192_ (.A(_089_),
    .Y(_093_));
 sky130_fd_sc_hd__nand2b_1 _193_ (.A_N(net19),
    .B(net18),
    .Y(_000_));
 sky130_fd_sc_hd__o31a_1 _194_ (.A1(net8),
    .A2(net6),
    .A3(net7),
    .B1(_000_),
    .X(_001_));
 sky130_fd_sc_hd__xnor2_1 _195_ (.A(net9),
    .B(_001_),
    .Y(_002_));
 sky130_fd_sc_hd__or2_1 _196_ (.A(net5),
    .B(_002_),
    .X(_003_));
 sky130_fd_sc_hd__o21a_1 _197_ (.A1(net6),
    .A2(net7),
    .B1(_000_),
    .X(_004_));
 sky130_fd_sc_hd__xnor2_1 _198_ (.A(net8),
    .B(_004_),
    .Y(_005_));
 sky130_fd_sc_hd__or2_1 _199_ (.A(net4),
    .B(_005_),
    .X(_006_));
 sky130_fd_sc_hd__nand3b_1 _200_ (.A_N(net7),
    .B(_000_),
    .C(net6),
    .Y(_007_));
 sky130_fd_sc_hd__a21bo_1 _201_ (.A1(net6),
    .A2(_000_),
    .B1_N(net7),
    .X(_008_));
 sky130_fd_sc_hd__a21o_1 _202_ (.A1(_007_),
    .A2(_008_),
    .B1(net3),
    .X(_009_));
 sky130_fd_sc_hd__or2b_1 _203_ (.A(net2),
    .B_N(net6),
    .X(_010_));
 sky130_fd_sc_hd__and3_1 _204_ (.A(net3),
    .B(_007_),
    .C(_008_),
    .X(_011_));
 sky130_fd_sc_hd__a21o_1 _205_ (.A1(_009_),
    .A2(_010_),
    .B1(_011_),
    .X(_012_));
 sky130_fd_sc_hd__and2_1 _206_ (.A(net5),
    .B(_002_),
    .X(_013_));
 sky130_fd_sc_hd__and2_1 _207_ (.A(net4),
    .B(_005_),
    .X(_014_));
 sky130_fd_sc_hd__a211o_1 _208_ (.A1(_006_),
    .A2(_012_),
    .B1(_013_),
    .C1(_014_),
    .X(_015_));
 sky130_fd_sc_hd__a21oi_1 _209_ (.A1(net9),
    .A2(_000_),
    .B1(_001_),
    .Y(_016_));
 sky130_fd_sc_hd__a21oi_1 _210_ (.A1(_003_),
    .A2(_015_),
    .B1(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__a31o_1 _211_ (.A1(_016_),
    .A2(_003_),
    .A3(_015_),
    .B1(net19),
    .X(_018_));
 sky130_fd_sc_hd__or2_1 _212_ (.A(_017_),
    .B(_018_),
    .X(_019_));
 sky130_fd_sc_hd__nand2b_1 _213_ (.A_N(net21),
    .B(net20),
    .Y(_020_));
 sky130_fd_sc_hd__o31a_1 _214_ (.A1(net16),
    .A2(net14),
    .A3(net15),
    .B1(_020_),
    .X(_021_));
 sky130_fd_sc_hd__xnor2_1 _215_ (.A(net17),
    .B(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__or2_1 _216_ (.A(net13),
    .B(_022_),
    .X(_023_));
 sky130_fd_sc_hd__o21a_1 _217_ (.A1(net14),
    .A2(net15),
    .B1(_020_),
    .X(_024_));
 sky130_fd_sc_hd__xnor2_1 _218_ (.A(net16),
    .B(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__or2_1 _219_ (.A(net12),
    .B(_025_),
    .X(_026_));
 sky130_fd_sc_hd__nand3b_1 _220_ (.A_N(net15),
    .B(_020_),
    .C(net14),
    .Y(_027_));
 sky130_fd_sc_hd__a21bo_1 _221_ (.A1(net14),
    .A2(_020_),
    .B1_N(net15),
    .X(_028_));
 sky130_fd_sc_hd__a21o_1 _222_ (.A1(_027_),
    .A2(_028_),
    .B1(net11),
    .X(_029_));
 sky130_fd_sc_hd__or2b_1 _223_ (.A(net10),
    .B_N(net14),
    .X(_030_));
 sky130_fd_sc_hd__and3_1 _224_ (.A(net11),
    .B(_027_),
    .C(_028_),
    .X(_031_));
 sky130_fd_sc_hd__a21o_1 _225_ (.A1(_029_),
    .A2(_030_),
    .B1(_031_),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _226_ (.A(net13),
    .B(_022_),
    .X(_033_));
 sky130_fd_sc_hd__and2_1 _227_ (.A(net12),
    .B(_025_),
    .X(_034_));
 sky130_fd_sc_hd__a211o_1 _228_ (.A1(_026_),
    .A2(_032_),
    .B1(_033_),
    .C1(_034_),
    .X(_035_));
 sky130_fd_sc_hd__a21oi_1 _229_ (.A1(net17),
    .A2(_020_),
    .B1(_021_),
    .Y(_036_));
 sky130_fd_sc_hd__a21oi_1 _230_ (.A1(_023_),
    .A2(_035_),
    .B1(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__a31o_1 _231_ (.A1(_036_),
    .A2(_023_),
    .A3(_035_),
    .B1(net21),
    .X(_038_));
 sky130_fd_sc_hd__or2_1 _232_ (.A(_037_),
    .B(_038_),
    .X(_039_));
 sky130_fd_sc_hd__nor3_2 _233_ (.A(_124_),
    .B(_037_),
    .C(_038_),
    .Y(net31));
 sky130_fd_sc_hd__nor3_1 _234_ (.A(_124_),
    .B(_017_),
    .C(_018_),
    .Y(net32));
 sky130_fd_sc_hd__o22a_1 _235_ (.A1(_019_),
    .A2(_039_),
    .B1(net31),
    .B2(net32),
    .X(net22));
 sky130_fd_sc_hd__inv_2 _236_ (.A(net19),
    .Y(_040_));
 sky130_fd_sc_hd__o2bb2a_1 _237_ (.A1_N(net6),
    .A2_N(net2),
    .B1(_040_),
    .B2(net18),
    .X(_041_));
 sky130_fd_sc_hd__o21a_1 _238_ (.A1(net6),
    .A2(net2),
    .B1(_041_),
    .X(_042_));
 sky130_fd_sc_hd__a31o_1 _239_ (.A1(net6),
    .A2(net19),
    .A3(net2),
    .B1(_042_),
    .X(_043_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(net21),
    .Y(_044_));
 sky130_fd_sc_hd__o2bb2a_1 _241_ (.A1_N(net14),
    .A2_N(net10),
    .B1(_044_),
    .B2(net20),
    .X(_045_));
 sky130_fd_sc_hd__o21a_1 _242_ (.A1(net14),
    .A2(net10),
    .B1(_045_),
    .X(_046_));
 sky130_fd_sc_hd__a31o_1 _243_ (.A1(net14),
    .A2(net21),
    .A3(net10),
    .B1(_046_),
    .X(_047_));
 sky130_fd_sc_hd__and2_1 _244_ (.A(_089_),
    .B(_047_),
    .X(_048_));
 sky130_fd_sc_hd__clkbuf_1 _245_ (.A(_048_),
    .X(net23));
 sky130_fd_sc_hd__and2_1 _246_ (.A(_089_),
    .B(_043_),
    .X(_049_));
 sky130_fd_sc_hd__clkbuf_1 _247_ (.A(_049_),
    .X(net27));
 sky130_fd_sc_hd__o2bb2a_1 _248_ (.A1_N(_043_),
    .A2_N(_047_),
    .B1(net23),
    .B2(net27),
    .X(net33));
 sky130_fd_sc_hd__or2b_1 _249_ (.A(_011_),
    .B_N(_009_),
    .X(_050_));
 sky130_fd_sc_hd__xnor2_1 _250_ (.A(_050_),
    .B(_010_),
    .Y(_051_));
 sky130_fd_sc_hd__o21a_1 _251_ (.A1(net7),
    .A2(net18),
    .B1(net3),
    .X(_052_));
 sky130_fd_sc_hd__a211o_1 _252_ (.A1(net7),
    .A2(net18),
    .B1(_040_),
    .C1(_052_),
    .X(_053_));
 sky130_fd_sc_hd__o21a_1 _253_ (.A1(net19),
    .A2(_051_),
    .B1(_053_),
    .X(_054_));
 sky130_fd_sc_hd__or2b_1 _254_ (.A(_031_),
    .B_N(_029_),
    .X(_055_));
 sky130_fd_sc_hd__xnor2_1 _255_ (.A(_055_),
    .B(_030_),
    .Y(_056_));
 sky130_fd_sc_hd__o21a_1 _256_ (.A1(net15),
    .A2(net20),
    .B1(net11),
    .X(_057_));
 sky130_fd_sc_hd__a211o_1 _257_ (.A1(net15),
    .A2(net20),
    .B1(_044_),
    .C1(_057_),
    .X(_058_));
 sky130_fd_sc_hd__o21a_1 _258_ (.A1(net21),
    .A2(_056_),
    .B1(_058_),
    .X(_059_));
 sky130_fd_sc_hd__and2_1 _259_ (.A(_089_),
    .B(_059_),
    .X(_060_));
 sky130_fd_sc_hd__clkbuf_1 _260_ (.A(_060_),
    .X(net24));
 sky130_fd_sc_hd__and2_1 _261_ (.A(_089_),
    .B(_054_),
    .X(_061_));
 sky130_fd_sc_hd__clkbuf_1 _262_ (.A(_061_),
    .X(net28));
 sky130_fd_sc_hd__o2bb2a_1 _263_ (.A1_N(_054_),
    .A2_N(_059_),
    .B1(net24),
    .B2(net28),
    .X(net34));
 sky130_fd_sc_hd__a21o_1 _264_ (.A1(net18),
    .A2(net4),
    .B1(net8),
    .X(_062_));
 sky130_fd_sc_hd__or2_1 _265_ (.A(net18),
    .B(net4),
    .X(_063_));
 sky130_fd_sc_hd__xor2_1 _266_ (.A(net4),
    .B(_005_),
    .X(_064_));
 sky130_fd_sc_hd__or2_1 _267_ (.A(_064_),
    .B(_012_),
    .X(_065_));
 sky130_fd_sc_hd__a21oi_1 _268_ (.A1(_064_),
    .A2(_012_),
    .B1(net19),
    .Y(_066_));
 sky130_fd_sc_hd__a32o_1 _269_ (.A1(net19),
    .A2(_062_),
    .A3(_063_),
    .B1(_065_),
    .B2(_066_),
    .X(_067_));
 sky130_fd_sc_hd__a21o_1 _270_ (.A1(net20),
    .A2(net12),
    .B1(net16),
    .X(_068_));
 sky130_fd_sc_hd__or2_1 _271_ (.A(net20),
    .B(net12),
    .X(_069_));
 sky130_fd_sc_hd__xor2_1 _272_ (.A(net12),
    .B(_025_),
    .X(_070_));
 sky130_fd_sc_hd__or2_1 _273_ (.A(_070_),
    .B(_032_),
    .X(_071_));
 sky130_fd_sc_hd__a21oi_1 _274_ (.A1(_070_),
    .A2(_032_),
    .B1(net21),
    .Y(_072_));
 sky130_fd_sc_hd__a32o_1 _275_ (.A1(net21),
    .A2(_068_),
    .A3(_069_),
    .B1(_071_),
    .B2(_072_),
    .X(_073_));
 sky130_fd_sc_hd__and2_1 _276_ (.A(net1),
    .B(_073_),
    .X(_074_));
 sky130_fd_sc_hd__clkbuf_1 _277_ (.A(_074_),
    .X(net25));
 sky130_fd_sc_hd__and2_1 _278_ (.A(_089_),
    .B(_067_),
    .X(_075_));
 sky130_fd_sc_hd__clkbuf_1 _279_ (.A(_075_),
    .X(net29));
 sky130_fd_sc_hd__o2bb2a_1 _280_ (.A1_N(_067_),
    .A2_N(_073_),
    .B1(net25),
    .B2(net29),
    .X(net35));
 sky130_fd_sc_hd__a21oi_1 _281_ (.A1(_006_),
    .A2(_012_),
    .B1(_014_),
    .Y(_076_));
 sky130_fd_sc_hd__and2b_1 _282_ (.A_N(_013_),
    .B(_003_),
    .X(_077_));
 sky130_fd_sc_hd__xnor2_1 _283_ (.A(_076_),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__nor2_1 _284_ (.A(net19),
    .B(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__o21a_1 _285_ (.A1(net9),
    .A2(net18),
    .B1(net5),
    .X(_080_));
 sky130_fd_sc_hd__a21o_1 _286_ (.A1(net9),
    .A2(net18),
    .B1(_040_),
    .X(_081_));
 sky130_fd_sc_hd__nor2_1 _287_ (.A(_080_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__a21o_1 _288_ (.A1(_026_),
    .A2(_032_),
    .B1(_034_),
    .X(_083_));
 sky130_fd_sc_hd__and2b_1 _289_ (.A_N(_033_),
    .B(_023_),
    .X(_084_));
 sky130_fd_sc_hd__xnor2_1 _290_ (.A(_083_),
    .B(_084_),
    .Y(_085_));
 sky130_fd_sc_hd__o21a_1 _291_ (.A1(net17),
    .A2(net20),
    .B1(net13),
    .X(_086_));
 sky130_fd_sc_hd__a211oi_2 _292_ (.A1(net17),
    .A2(net20),
    .B1(_044_),
    .C1(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__a21o_1 _293_ (.A1(_044_),
    .A2(_085_),
    .B1(_087_),
    .X(_088_));
 sky130_fd_sc_hd__a211oi_2 _294_ (.A1(_044_),
    .A2(_085_),
    .B1(_087_),
    .C1(_124_),
    .Y(net26));
 sky130_fd_sc_hd__o221a_1 _295_ (.A1(net19),
    .A2(_078_),
    .B1(_080_),
    .B2(_081_),
    .C1(_089_),
    .X(net30));
 sky130_fd_sc_hd__o32a_1 _296_ (.A1(_079_),
    .A2(_082_),
    .A3(_088_),
    .B1(net26),
    .B2(net30),
    .X(net36));
 sky130_fd_sc_hd__conb_1 macro_decap_12_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 macro_decap_12_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 macro_decap_12_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 macro_decap_12_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 macro_decap_12_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 macro_decap_12_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 macro_decap_12_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 macro_decap_12_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 macro_decap_12_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 macro_decap_12_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 macro_decap_12_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 macro_decap_12_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 macro_decap_12_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 macro_decap_12_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 macro_decap_12_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 macro_decap_12_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 macro_decap_12_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 macro_decap_12_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 macro_decap_12_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 macro_decap_12_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 macro_decap_12_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 macro_decap_12_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 macro_decap_12_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 macro_decap_12_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 macro_decap_12_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 macro_decap_12_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 macro_decap_12_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 macro_decap_12_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 macro_decap_12_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 macro_decap_12_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 macro_decap_12_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 macro_decap_12_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 macro_decap_12_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 macro_decap_12_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 macro_decap_12_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 macro_decap_12_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 macro_decap_12_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 macro_decap_12_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 macro_decap_12_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 macro_decap_12_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 macro_decap_12_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 macro_decap_12_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 macro_decap_12_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 macro_decap_12_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 macro_decap_12_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 macro_decap_12_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 macro_decap_12_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 macro_decap_12_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 macro_decap_12_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 macro_decap_12_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 macro_decap_12_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 macro_decap_12_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 macro_decap_12_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 macro_decap_12_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 macro_decap_12_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 macro_decap_12_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 macro_decap_12_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 macro_decap_12_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 macro_decap_12_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 macro_decap_12_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 macro_decap_12_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 macro_decap_12_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 macro_decap_12_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 macro_decap_12_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 macro_decap_12_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 macro_decap_12_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 macro_decap_12_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 macro_decap_12_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 macro_decap_12_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 macro_decap_12_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 macro_decap_12_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 macro_decap_12_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 macro_decap_12_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 macro_decap_12_111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 macro_decap_12_112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 macro_decap_12_113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 macro_decap_12_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 macro_decap_12_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 macro_decap_12_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 macro_decap_12_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 macro_decap_12_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 macro_decap_12_119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 macro_decap_12_120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 macro_decap_12_121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 macro_decap_12_122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 macro_decap_12_123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 macro_decap_12_124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 macro_decap_12_125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 macro_decap_12_126 (.LO(net126));
 sky130_fd_sc_hd__conb_1 macro_decap_12_127 (.LO(net127));
 sky130_fd_sc_hd__conb_1 macro_decap_12_128 (.LO(net128));
 sky130_fd_sc_hd__conb_1 macro_decap_12_129 (.LO(net129));
 sky130_fd_sc_hd__conb_1 macro_decap_12_130 (.LO(net130));
 sky130_fd_sc_hd__conb_1 macro_decap_12_131 (.LO(net131));
 sky130_fd_sc_hd__conb_1 macro_decap_12_132 (.LO(net132));
 sky130_fd_sc_hd__conb_1 macro_decap_12_133 (.LO(net133));
 sky130_fd_sc_hd__conb_1 macro_decap_12_134 (.LO(net134));
 sky130_fd_sc_hd__conb_1 macro_decap_12_135 (.LO(net135));
 sky130_fd_sc_hd__conb_1 macro_decap_12_136 (.LO(net136));
 sky130_fd_sc_hd__conb_1 macro_decap_12_137 (.LO(net137));
 sky130_fd_sc_hd__conb_1 macro_decap_12_138 (.LO(net138));
 sky130_fd_sc_hd__conb_1 macro_decap_12_139 (.LO(net139));
 sky130_fd_sc_hd__conb_1 macro_decap_12_140 (.LO(net140));
 sky130_fd_sc_hd__conb_1 macro_decap_12_141 (.LO(net141));
 sky130_fd_sc_hd__conb_1 macro_decap_12_142 (.LO(net142));
 sky130_fd_sc_hd__conb_1 macro_decap_12_143 (.LO(net143));
 sky130_fd_sc_hd__conb_1 macro_decap_12_144 (.LO(net144));
 sky130_fd_sc_hd__conb_1 macro_decap_12_145 (.LO(net145));
 sky130_fd_sc_hd__conb_1 macro_decap_12_146 (.LO(net146));
 sky130_fd_sc_hd__conb_1 macro_decap_12_147 (.LO(net147));
 sky130_fd_sc_hd__conb_1 macro_decap_12_148 (.LO(net148));
 sky130_fd_sc_hd__conb_1 macro_decap_12_149 (.LO(net149));
 sky130_fd_sc_hd__conb_1 macro_decap_12_150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 macro_decap_12_151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 macro_decap_12_152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 macro_decap_12_153 (.LO(net153));
 sky130_fd_sc_hd__conb_1 macro_decap_12_154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 macro_decap_12_155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 macro_decap_12_156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 macro_decap_12_157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 macro_decap_12_158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 macro_decap_12_159 (.LO(net159));
 sky130_fd_sc_hd__conb_1 macro_decap_12_160 (.LO(net160));
 sky130_fd_sc_hd__conb_1 macro_decap_12_161 (.LO(net161));
 sky130_fd_sc_hd__conb_1 macro_decap_12_162 (.LO(net162));
 sky130_fd_sc_hd__conb_1 macro_decap_12_163 (.LO(net163));
 sky130_fd_sc_hd__conb_1 macro_decap_12_164 (.LO(net164));
 sky130_fd_sc_hd__conb_1 macro_decap_12_165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 macro_decap_12_166 (.LO(net166));
 sky130_fd_sc_hd__conb_1 macro_decap_12_167 (.LO(net167));
 sky130_fd_sc_hd__conb_1 macro_decap_12_168 (.LO(net168));
 sky130_fd_sc_hd__conb_1 macro_decap_12_169 (.LO(net169));
 sky130_fd_sc_hd__conb_1 macro_decap_12_170 (.LO(net170));
 sky130_fd_sc_hd__conb_1 macro_decap_12_171 (.LO(net171));
 sky130_fd_sc_hd__conb_1 macro_decap_12_172 (.LO(net172));
 sky130_fd_sc_hd__conb_1 macro_decap_12_173 (.LO(net173));
 sky130_fd_sc_hd__conb_1 macro_decap_12_174 (.LO(net174));
 sky130_fd_sc_hd__conb_1 macro_decap_12_175 (.LO(net175));
 sky130_fd_sc_hd__conb_1 macro_decap_12_176 (.LO(net176));
 sky130_fd_sc_hd__conb_1 macro_decap_12_177 (.LO(net177));
 sky130_fd_sc_hd__conb_1 macro_decap_12_178 (.LO(net178));
 sky130_fd_sc_hd__conb_1 macro_decap_12_179 (.LO(net179));
 sky130_fd_sc_hd__conb_1 macro_decap_12_180 (.LO(net180));
 sky130_fd_sc_hd__conb_1 macro_decap_12_181 (.LO(net181));
 sky130_fd_sc_hd__conb_1 macro_decap_12_182 (.LO(net182));
 sky130_fd_sc_hd__conb_1 macro_decap_12_183 (.LO(net183));
 sky130_fd_sc_hd__conb_1 macro_decap_12_184 (.LO(net184));
 sky130_fd_sc_hd__conb_1 macro_decap_12_185 (.LO(net185));
 sky130_fd_sc_hd__conb_1 macro_decap_12_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 macro_decap_12_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 macro_decap_12_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 macro_decap_12_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 macro_decap_12_190 (.LO(net190));
 sky130_fd_sc_hd__conb_1 macro_decap_12_191 (.LO(net191));
 sky130_fd_sc_hd__conb_1 macro_decap_12_192 (.LO(net192));
 sky130_fd_sc_hd__conb_1 macro_decap_12_193 (.LO(net193));
 sky130_fd_sc_hd__conb_1 _519__194 (.LO(net194));
 sky130_fd_sc_hd__conb_1 _520__195 (.LO(net195));
 sky130_fd_sc_hd__conb_1 _521__196 (.LO(net196));
 sky130_fd_sc_hd__conb_1 _522__197 (.LO(net197));
 sky130_fd_sc_hd__conb_1 _523__198 (.LO(net198));
 sky130_fd_sc_hd__conb_1 _524__199 (.LO(net199));
 sky130_fd_sc_hd__conb_1 _525__200 (.LO(net200));
 sky130_fd_sc_hd__conb_1 _526__201 (.LO(net201));
 sky130_fd_sc_hd__conb_1 _527__202 (.LO(net202));
 sky130_fd_sc_hd__conb_1 _528__203 (.LO(net203));
 sky130_fd_sc_hd__conb_1 _529__204 (.LO(net204));
 sky130_fd_sc_hd__conb_1 _530__205 (.LO(net205));
 sky130_fd_sc_hd__conb_1 _531__206 (.LO(net206));
 sky130_fd_sc_hd__conb_1 _532__207 (.LO(net207));
 sky130_fd_sc_hd__conb_1 _533__208 (.LO(net208));
 sky130_fd_sc_hd__conb_1 _534__209 (.LO(net209));
 sky130_fd_sc_hd__conb_1 _535__210 (.LO(net210));
 sky130_fd_sc_hd__conb_1 _536__211 (.LO(net211));
 sky130_fd_sc_hd__conb_1 _537__212 (.LO(net212));
 sky130_fd_sc_hd__conb_1 _538__213 (.LO(net213));
 sky130_fd_sc_hd__conb_1 _539__214 (.LO(net214));
 sky130_fd_sc_hd__conb_1 _540__215 (.LO(net215));
 sky130_fd_sc_hd__conb_1 _541__216 (.LO(net216));
 sky130_fd_sc_hd__conb_1 _542__217 (.LO(net217));
 sky130_fd_sc_hd__conb_1 _543__218 (.LO(net218));
 sky130_fd_sc_hd__conb_1 _544__219 (.LO(net219));
 sky130_fd_sc_hd__conb_1 _545__220 (.LO(net220));
 sky130_fd_sc_hd__conb_1 _546__221 (.LO(net221));
 sky130_fd_sc_hd__conb_1 _547__222 (.LO(net222));
 sky130_fd_sc_hd__conb_1 _548__223 (.LO(net223));
 sky130_fd_sc_hd__conb_1 _549__224 (.LO(net224));
 sky130_fd_sc_hd__conb_1 _550__225 (.LO(net225));
 sky130_fd_sc_hd__conb_1 macro_decap_12_226 (.LO(net226));
 sky130_fd_sc_hd__conb_1 macro_decap_12_227 (.LO(net227));
 sky130_fd_sc_hd__conb_1 macro_decap_12_228 (.LO(net228));
 sky130_fd_sc_hd__conb_1 macro_decap_12_229 (.LO(net229));
 sky130_fd_sc_hd__conb_1 macro_decap_12_230 (.LO(net230));
 sky130_fd_sc_hd__conb_1 macro_decap_12_231 (.LO(net231));
 sky130_fd_sc_hd__conb_1 macro_decap_12_232 (.LO(net232));
 sky130_fd_sc_hd__conb_1 macro_decap_12_233 (.LO(net233));
 sky130_fd_sc_hd__conb_1 macro_decap_12_234 (.LO(net234));
 sky130_fd_sc_hd__conb_1 macro_decap_12_235 (.LO(net235));
 sky130_fd_sc_hd__conb_1 macro_decap_12_236 (.LO(net236));
 sky130_fd_sc_hd__conb_1 macro_decap_12_237 (.LO(net237));
 sky130_fd_sc_hd__conb_1 macro_decap_12_238 (.LO(net238));
 sky130_fd_sc_hd__conb_1 macro_decap_12_239 (.LO(net239));
 sky130_fd_sc_hd__conb_1 macro_decap_12_240 (.LO(net240));
 sky130_fd_sc_hd__conb_1 macro_decap_12_241 (.LO(net241));
 sky130_fd_sc_hd__conb_1 macro_decap_12_242 (.LO(net242));
 sky130_fd_sc_hd__conb_1 macro_decap_12_243 (.LO(net243));
 sky130_fd_sc_hd__conb_1 macro_decap_12_244 (.LO(net244));
 sky130_fd_sc_hd__conb_1 macro_decap_12_245 (.LO(net245));
 sky130_fd_sc_hd__conb_1 macro_decap_12_246 (.LO(net246));
 sky130_fd_sc_hd__conb_1 macro_decap_12_247 (.LO(net247));
 sky130_fd_sc_hd__conb_1 macro_decap_12_248 (.LO(net248));
 sky130_fd_sc_hd__conb_1 macro_decap_12_249 (.LO(net249));
 sky130_fd_sc_hd__conb_1 macro_decap_12_250 (.LO(net250));
 sky130_fd_sc_hd__conb_1 macro_decap_12_251 (.LO(net251));
 sky130_fd_sc_hd__conb_1 macro_decap_12_252 (.LO(net252));
 sky130_fd_sc_hd__conb_1 macro_decap_12_253 (.LO(net253));
 sky130_fd_sc_hd__conb_1 macro_decap_12_254 (.LO(net254));
 sky130_fd_sc_hd__conb_1 macro_decap_12_255 (.LO(net255));
 sky130_fd_sc_hd__conb_1 macro_decap_12_256 (.LO(net256));
 sky130_fd_sc_hd__conb_1 macro_decap_12_257 (.LO(net257));
 sky130_fd_sc_hd__conb_1 macro_decap_12_258 (.LO(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__C1 (.DIODE(_089_));
 sky130_fd_sc_hd__ebufn_8 _519_ (.A(net194),
    .TE_B(_093_),
    .Z(la_data_out[32]));
 sky130_fd_sc_hd__ebufn_8 _520_ (.A(net195),
    .TE_B(_094_),
    .Z(la_data_out[33]));
 sky130_fd_sc_hd__ebufn_8 _521_ (.A(net196),
    .TE_B(_095_),
    .Z(la_data_out[34]));
 sky130_fd_sc_hd__ebufn_8 _522_ (.A(net197),
    .TE_B(_096_),
    .Z(la_data_out[35]));
 sky130_fd_sc_hd__ebufn_8 _523_ (.A(net198),
    .TE_B(_097_),
    .Z(la_data_out[36]));
 sky130_fd_sc_hd__ebufn_8 _524_ (.A(net199),
    .TE_B(_098_),
    .Z(la_data_out[37]));
 sky130_fd_sc_hd__ebufn_8 _525_ (.A(net200),
    .TE_B(_099_),
    .Z(la_data_out[38]));
 sky130_fd_sc_hd__ebufn_8 _526_ (.A(net201),
    .TE_B(_100_),
    .Z(la_data_out[39]));
 sky130_fd_sc_hd__ebufn_8 _527_ (.A(net202),
    .TE_B(_101_),
    .Z(la_data_out[40]));
 sky130_fd_sc_hd__ebufn_8 _528_ (.A(net203),
    .TE_B(_102_),
    .Z(la_data_out[41]));
 sky130_fd_sc_hd__ebufn_8 _529_ (.A(net204),
    .TE_B(_103_),
    .Z(la_data_out[42]));
 sky130_fd_sc_hd__ebufn_8 _530_ (.A(net205),
    .TE_B(_104_),
    .Z(la_data_out[43]));
 sky130_fd_sc_hd__ebufn_8 _531_ (.A(net206),
    .TE_B(_105_),
    .Z(la_data_out[44]));
 sky130_fd_sc_hd__ebufn_8 _532_ (.A(net207),
    .TE_B(_106_),
    .Z(la_data_out[45]));
 sky130_fd_sc_hd__ebufn_8 _533_ (.A(net208),
    .TE_B(_107_),
    .Z(la_data_out[46]));
 sky130_fd_sc_hd__ebufn_8 _534_ (.A(net209),
    .TE_B(_108_),
    .Z(la_data_out[47]));
 sky130_fd_sc_hd__ebufn_8 _535_ (.A(net210),
    .TE_B(_109_),
    .Z(la_data_out[48]));
 sky130_fd_sc_hd__ebufn_8 _536_ (.A(net211),
    .TE_B(_110_),
    .Z(la_data_out[49]));
 sky130_fd_sc_hd__ebufn_8 _537_ (.A(net212),
    .TE_B(_111_),
    .Z(la_data_out[50]));
 sky130_fd_sc_hd__ebufn_8 _538_ (.A(net213),
    .TE_B(_112_),
    .Z(la_data_out[51]));
 sky130_fd_sc_hd__ebufn_8 _539_ (.A(net214),
    .TE_B(_113_),
    .Z(la_data_out[52]));
 sky130_fd_sc_hd__ebufn_8 _540_ (.A(net215),
    .TE_B(_114_),
    .Z(la_data_out[53]));
 sky130_fd_sc_hd__ebufn_8 _541_ (.A(net216),
    .TE_B(_115_),
    .Z(la_data_out[54]));
 sky130_fd_sc_hd__ebufn_8 _542_ (.A(net217),
    .TE_B(_116_),
    .Z(la_data_out[55]));
 sky130_fd_sc_hd__ebufn_8 _543_ (.A(net218),
    .TE_B(_117_),
    .Z(la_data_out[56]));
 sky130_fd_sc_hd__ebufn_8 _544_ (.A(net219),
    .TE_B(_118_),
    .Z(la_data_out[57]));
 sky130_fd_sc_hd__ebufn_8 _545_ (.A(net220),
    .TE_B(_119_),
    .Z(la_data_out[58]));
 sky130_fd_sc_hd__ebufn_8 _546_ (.A(net221),
    .TE_B(_120_),
    .Z(la_data_out[59]));
 sky130_fd_sc_hd__ebufn_8 _547_ (.A(net222),
    .TE_B(_121_),
    .Z(la_data_out[60]));
 sky130_fd_sc_hd__ebufn_8 _548_ (.A(net223),
    .TE_B(_122_),
    .Z(la_data_out[61]));
 sky130_fd_sc_hd__ebufn_8 _549_ (.A(net224),
    .TE_B(_123_),
    .Z(la_data_out[62]));
 sky130_fd_sc_hd__ebufn_8 _550_ (.A(net225),
    .TE_B(_124_),
    .Z(la_data_out[63]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_active),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[18]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[19]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(io_in[20]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[21]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[22]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(io_in[23]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(io_in[24]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(io_in[25]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(io_in[26]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(io_in[27]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(io_in[28]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(io_in[29]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(io_in[30]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(io_in[31]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(io_in[32]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(io_in[33]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(io_in[34]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(io_in[35]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(io_in[36]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(io_in[37]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(io_out[9]));
 sky130_fd_sc_hd__conb_1 macro_decap_12_37 (.LO(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__278__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__261__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__259__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__246__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__170__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__159__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_active));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(io_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(io_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(io_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__157__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__286__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__285__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__265__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__284__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__269__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__253__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__236__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__A_N (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__274__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__231__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__A_N (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__B1 (.DIODE(net31));
 sky130_fd_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_580 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_566 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_578 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_590 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_150 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_547 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_554 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_416 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_420 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_444 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_384 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_384 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_396 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_408 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_348 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_356 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_328 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_322 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_329 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_311 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_38_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_40_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_42_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_44_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_46_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_48_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_50_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_52_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_54_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_56_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_58_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_60_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_62_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_64_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_66_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_68_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_70_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_72_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_74_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_76_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_78_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_80_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_82_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_84_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_86_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_88_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_349 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_361 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_321 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_90_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_305 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_357 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_380 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_405 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_265 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_277 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_333 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_339 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_377 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_389 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_433 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_445 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_92_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_293 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_358 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_364 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_388 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_417 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_423 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_473 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_373 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_379 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_391 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_443 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_450 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_94_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_237 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_249 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_461 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_469 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_221 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_489 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_501 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_96_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_486 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_492 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_517 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_573 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_585 ();
 sky130_fd_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_41 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_109 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_153 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_165 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_209 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_456 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_492 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_498 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_545 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_557 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_601 ();
 sky130_fd_sc_hd__decap_12 FILLER_98_613 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_69 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_81 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_413 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_529 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_565 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_577 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_589 ();
 sky130_fd_sc_hd__decap_12 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_143 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_173 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_400 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_594 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_600 ();
 sky130_fd_sc_hd__decap_12 FILLER_100_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_624 ();
 sky130_fd_sc_hd__decap_12 FILLER_101_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_57 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_617 ();
 assign io_oeb[0] = net226;
 assign io_oeb[10] = net236;
 assign io_oeb[11] = net237;
 assign io_oeb[12] = net238;
 assign io_oeb[13] = net239;
 assign io_oeb[14] = net240;
 assign io_oeb[15] = net241;
 assign io_oeb[16] = net242;
 assign io_oeb[17] = net243;
 assign io_oeb[18] = net244;
 assign io_oeb[19] = net245;
 assign io_oeb[1] = net227;
 assign io_oeb[20] = net246;
 assign io_oeb[21] = net247;
 assign io_oeb[22] = net248;
 assign io_oeb[23] = net249;
 assign io_oeb[24] = net250;
 assign io_oeb[25] = net251;
 assign io_oeb[26] = net252;
 assign io_oeb[27] = net253;
 assign io_oeb[28] = net254;
 assign io_oeb[29] = net255;
 assign io_oeb[2] = net228;
 assign io_oeb[30] = net256;
 assign io_oeb[31] = net257;
 assign io_oeb[32] = net258;
 assign io_oeb[33] = net37;
 assign io_oeb[34] = net38;
 assign io_oeb[35] = net39;
 assign io_oeb[36] = net40;
 assign io_oeb[37] = net41;
 assign io_oeb[3] = net229;
 assign io_oeb[4] = net230;
 assign io_oeb[5] = net231;
 assign io_oeb[6] = net232;
 assign io_oeb[7] = net233;
 assign io_oeb[8] = net234;
 assign io_oeb[9] = net235;
 assign io_out[18] = net45;
 assign io_out[19] = net46;
 assign io_out[1] = net42;
 assign io_out[20] = net47;
 assign io_out[21] = net48;
 assign io_out[22] = net49;
 assign io_out[23] = net50;
 assign io_out[24] = net51;
 assign io_out[25] = net52;
 assign io_out[26] = net53;
 assign io_out[27] = net54;
 assign io_out[28] = net55;
 assign io_out[29] = net56;
 assign io_out[2] = net43;
 assign io_out[30] = net57;
 assign io_out[31] = net58;
 assign io_out[32] = net59;
 assign io_out[33] = net60;
 assign io_out[34] = net61;
 assign io_out[35] = net62;
 assign io_out[36] = net63;
 assign io_out[37] = net64;
 assign io_out[3] = net44;
 assign la_data_out[0] = net65;
 assign la_data_out[100] = net133;
 assign la_data_out[101] = net134;
 assign la_data_out[102] = net135;
 assign la_data_out[103] = net136;
 assign la_data_out[104] = net137;
 assign la_data_out[105] = net138;
 assign la_data_out[106] = net139;
 assign la_data_out[107] = net140;
 assign la_data_out[108] = net141;
 assign la_data_out[109] = net142;
 assign la_data_out[10] = net75;
 assign la_data_out[110] = net143;
 assign la_data_out[111] = net144;
 assign la_data_out[112] = net145;
 assign la_data_out[113] = net146;
 assign la_data_out[114] = net147;
 assign la_data_out[115] = net148;
 assign la_data_out[116] = net149;
 assign la_data_out[117] = net150;
 assign la_data_out[118] = net151;
 assign la_data_out[119] = net152;
 assign la_data_out[11] = net76;
 assign la_data_out[120] = net153;
 assign la_data_out[121] = net154;
 assign la_data_out[122] = net155;
 assign la_data_out[123] = net156;
 assign la_data_out[124] = net157;
 assign la_data_out[125] = net158;
 assign la_data_out[126] = net159;
 assign la_data_out[127] = net160;
 assign la_data_out[12] = net77;
 assign la_data_out[13] = net78;
 assign la_data_out[14] = net79;
 assign la_data_out[15] = net80;
 assign la_data_out[16] = net81;
 assign la_data_out[17] = net82;
 assign la_data_out[18] = net83;
 assign la_data_out[19] = net84;
 assign la_data_out[1] = net66;
 assign la_data_out[20] = net85;
 assign la_data_out[21] = net86;
 assign la_data_out[22] = net87;
 assign la_data_out[23] = net88;
 assign la_data_out[24] = net89;
 assign la_data_out[25] = net90;
 assign la_data_out[26] = net91;
 assign la_data_out[27] = net92;
 assign la_data_out[28] = net93;
 assign la_data_out[29] = net94;
 assign la_data_out[2] = net67;
 assign la_data_out[30] = net95;
 assign la_data_out[31] = net96;
 assign la_data_out[3] = net68;
 assign la_data_out[4] = net69;
 assign la_data_out[5] = net70;
 assign la_data_out[64] = net97;
 assign la_data_out[65] = net98;
 assign la_data_out[66] = net99;
 assign la_data_out[67] = net100;
 assign la_data_out[68] = net101;
 assign la_data_out[69] = net102;
 assign la_data_out[6] = net71;
 assign la_data_out[70] = net103;
 assign la_data_out[71] = net104;
 assign la_data_out[72] = net105;
 assign la_data_out[73] = net106;
 assign la_data_out[74] = net107;
 assign la_data_out[75] = net108;
 assign la_data_out[76] = net109;
 assign la_data_out[77] = net110;
 assign la_data_out[78] = net111;
 assign la_data_out[79] = net112;
 assign la_data_out[7] = net72;
 assign la_data_out[80] = net113;
 assign la_data_out[81] = net114;
 assign la_data_out[82] = net115;
 assign la_data_out[83] = net116;
 assign la_data_out[84] = net117;
 assign la_data_out[85] = net118;
 assign la_data_out[86] = net119;
 assign la_data_out[87] = net120;
 assign la_data_out[88] = net121;
 assign la_data_out[89] = net122;
 assign la_data_out[8] = net73;
 assign la_data_out[90] = net123;
 assign la_data_out[91] = net124;
 assign la_data_out[92] = net125;
 assign la_data_out[93] = net126;
 assign la_data_out[94] = net127;
 assign la_data_out[95] = net128;
 assign la_data_out[96] = net129;
 assign la_data_out[97] = net130;
 assign la_data_out[98] = net131;
 assign la_data_out[99] = net132;
 assign la_data_out[9] = net74;
 assign wbs_ack_o = net161;
 assign wbs_dat_o[0] = net162;
 assign wbs_dat_o[10] = net172;
 assign wbs_dat_o[11] = net173;
 assign wbs_dat_o[12] = net174;
 assign wbs_dat_o[13] = net175;
 assign wbs_dat_o[14] = net176;
 assign wbs_dat_o[15] = net177;
 assign wbs_dat_o[16] = net178;
 assign wbs_dat_o[17] = net179;
 assign wbs_dat_o[18] = net180;
 assign wbs_dat_o[19] = net181;
 assign wbs_dat_o[1] = net163;
 assign wbs_dat_o[20] = net182;
 assign wbs_dat_o[21] = net183;
 assign wbs_dat_o[22] = net184;
 assign wbs_dat_o[23] = net185;
 assign wbs_dat_o[24] = net186;
 assign wbs_dat_o[25] = net187;
 assign wbs_dat_o[26] = net188;
 assign wbs_dat_o[27] = net189;
 assign wbs_dat_o[28] = net190;
 assign wbs_dat_o[29] = net191;
 assign wbs_dat_o[2] = net164;
 assign wbs_dat_o[30] = net192;
 assign wbs_dat_o[31] = net193;
 assign wbs_dat_o[3] = net165;
 assign wbs_dat_o[4] = net166;
 assign wbs_dat_o[5] = net167;
 assign wbs_dat_o[6] = net168;
 assign wbs_dat_o[7] = net169;
 assign wbs_dat_o[8] = net170;
 assign wbs_dat_o[9] = net171;
endmodule

