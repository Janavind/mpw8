magic
tech sky130A
magscale 1 2
timestamp 1672276709
<< viali >>
rect 5365 57545 5399 57579
rect 11161 57545 11195 57579
rect 12173 57545 12207 57579
rect 13553 57545 13587 57579
rect 15025 57545 15059 57579
rect 16957 57545 16991 57579
rect 17693 57545 17727 57579
rect 19073 57545 19107 57579
rect 20821 57545 20855 57579
rect 21833 57545 21867 57579
rect 23121 57545 23155 57579
rect 23949 57545 23983 57579
rect 40049 57545 40083 57579
rect 41981 57545 42015 57579
rect 48007 57545 48041 57579
rect 52653 57545 52687 57579
rect 3893 57477 3927 57511
rect 34713 57477 34747 57511
rect 52929 57477 52963 57511
rect 4537 57409 4571 57443
rect 5549 57409 5583 57443
rect 6469 57409 6503 57443
rect 7757 57409 7791 57443
rect 8585 57409 8619 57443
rect 9321 57409 9355 57443
rect 10241 57409 10275 57443
rect 11345 57409 11379 57443
rect 12357 57409 12391 57443
rect 13737 57409 13771 57443
rect 14197 57409 14231 57443
rect 15209 57409 15243 57443
rect 15761 57409 15795 57443
rect 17141 57409 17175 57443
rect 17877 57409 17911 57443
rect 19257 57409 19291 57443
rect 19901 57409 19935 57443
rect 21005 57409 21039 57443
rect 22017 57409 22051 57443
rect 23305 57409 23339 57443
rect 23765 57409 23799 57443
rect 24777 57409 24811 57443
rect 25605 57409 25639 57443
rect 26893 57409 26927 57443
rect 27169 57409 27203 57443
rect 27629 57409 27663 57443
rect 27905 57409 27939 57443
rect 29101 57409 29135 57443
rect 29285 57409 29319 57443
rect 29561 57409 29595 57443
rect 30389 57409 30423 57443
rect 31401 57409 31435 57443
rect 32321 57409 32355 57443
rect 37473 57409 37507 57443
rect 39497 57409 39531 57443
rect 40233 57409 40267 57443
rect 41245 57409 41279 57443
rect 41429 57409 41463 57443
rect 43361 57409 43395 57443
rect 44097 57409 44131 57443
rect 46029 57409 46063 57443
rect 46765 57409 46799 57443
rect 47777 57409 47811 57443
rect 49801 57409 49835 57443
rect 51641 57409 51675 57443
rect 53941 57409 53975 57443
rect 54677 57409 54711 57443
rect 55505 57409 55539 57443
rect 56241 57409 56275 57443
rect 24961 57341 24995 57375
rect 25789 57341 25823 57375
rect 29377 57341 29411 57375
rect 31677 57341 31711 57375
rect 32597 57341 32631 57375
rect 36185 57341 36219 57375
rect 36461 57341 36495 57375
rect 38117 57341 38151 57375
rect 38393 57341 38427 57375
rect 40325 57341 40359 57375
rect 40417 57341 40451 57375
rect 40509 57341 40543 57375
rect 43085 57341 43119 57375
rect 44373 57341 44407 57375
rect 50077 57341 50111 57375
rect 4077 57273 4111 57307
rect 27813 57273 27847 57307
rect 28917 57273 28951 57307
rect 29193 57273 29227 57307
rect 30573 57273 30607 57307
rect 49065 57273 49099 57307
rect 51825 57273 51859 57307
rect 7297 57205 7331 57239
rect 24593 57205 24627 57239
rect 25421 57205 25455 57239
rect 27721 57205 27755 57239
rect 31217 57205 31251 57239
rect 31585 57205 31619 57239
rect 33701 57205 33735 57239
rect 34805 57205 34839 57239
rect 35357 57205 35391 57239
rect 41061 57205 41095 57239
rect 43913 57205 43947 57239
rect 44281 57205 44315 57239
rect 44833 57205 44867 57239
rect 45937 57205 45971 57239
rect 46581 57205 46615 57239
rect 54125 57205 54159 57239
rect 55689 57205 55723 57239
rect 3709 57001 3743 57035
rect 6101 57001 6135 57035
rect 7481 57001 7515 57035
rect 11621 57001 11655 57035
rect 13001 57001 13035 57035
rect 17141 57001 17175 57035
rect 19165 57001 19199 57035
rect 21281 57001 21315 57035
rect 24317 57001 24351 57035
rect 25697 57001 25731 57035
rect 27169 57001 27203 57035
rect 28641 57001 28675 57035
rect 29929 57001 29963 57035
rect 31033 57001 31067 57035
rect 31677 57001 31711 57035
rect 34253 57001 34287 57035
rect 35173 57001 35207 57035
rect 43269 57001 43303 57035
rect 47501 57001 47535 57035
rect 49709 57001 49743 57035
rect 50813 57001 50847 57035
rect 52101 57001 52135 57035
rect 52745 57001 52779 57035
rect 53389 57001 53423 57035
rect 54033 57001 54067 57035
rect 54861 57001 54895 57035
rect 55505 57001 55539 57035
rect 56241 57001 56275 57035
rect 22385 56933 22419 56967
rect 27721 56933 27755 56967
rect 30481 56933 30515 56967
rect 32229 56933 32263 56967
rect 36093 56933 36127 56967
rect 46857 56933 46891 56967
rect 51457 56933 51491 56967
rect 12357 56865 12391 56899
rect 23673 56865 23707 56899
rect 25053 56865 25087 56899
rect 27077 56865 27111 56899
rect 29469 56865 29503 56899
rect 37841 56865 37875 56899
rect 38209 56865 38243 56899
rect 38945 56865 38979 56899
rect 40601 56865 40635 56899
rect 43913 56865 43947 56899
rect 48421 56865 48455 56899
rect 22569 56797 22603 56831
rect 23765 56797 23799 56831
rect 24192 56797 24226 56831
rect 25145 56797 25179 56831
rect 25572 56797 25606 56831
rect 26341 56797 26375 56831
rect 26433 56797 26467 56831
rect 27540 56797 27574 56831
rect 28365 56797 28399 56831
rect 28457 56797 28491 56831
rect 28733 56797 28767 56831
rect 29193 56797 29227 56831
rect 29377 56797 29411 56831
rect 29561 56797 29595 56831
rect 29745 56797 29779 56831
rect 31802 56797 31836 56831
rect 32321 56797 32355 56831
rect 33425 56797 33459 56831
rect 33517 56797 33551 56831
rect 33701 56797 33735 56831
rect 33793 56797 33827 56831
rect 35541 56797 35575 56831
rect 36001 56797 36035 56831
rect 36277 56797 36311 56831
rect 36553 56797 36587 56831
rect 36829 56797 36863 56831
rect 37381 56797 37415 56831
rect 38025 56797 38059 56831
rect 38117 56797 38151 56831
rect 38301 56797 38335 56831
rect 39221 56797 39255 56831
rect 40509 56797 40543 56831
rect 41028 56797 41062 56831
rect 41797 56797 41831 56831
rect 41889 56797 41923 56831
rect 42085 56797 42119 56831
rect 42175 56797 42209 56831
rect 42901 56797 42935 56831
rect 43085 56797 43119 56831
rect 43361 56797 43395 56831
rect 44097 56797 44131 56831
rect 44465 56797 44499 56831
rect 44741 56797 44775 56831
rect 45201 56797 45235 56831
rect 45845 56797 45879 56831
rect 48697 56797 48731 56831
rect 28181 56729 28215 56763
rect 35357 56729 35391 56763
rect 44005 56729 44039 56763
rect 23121 56661 23155 56695
rect 24133 56661 24167 56695
rect 25513 56661 25547 56695
rect 26157 56661 26191 56695
rect 27537 56661 27571 56695
rect 31861 56661 31895 56695
rect 33241 56661 33275 56695
rect 40969 56661 41003 56695
rect 41153 56661 41187 56695
rect 41613 56661 41647 56695
rect 23581 56457 23615 56491
rect 28457 56457 28491 56491
rect 32045 56457 32079 56491
rect 33977 56457 34011 56491
rect 35541 56457 35575 56491
rect 37013 56457 37047 56491
rect 39589 56457 39623 56491
rect 40969 56457 41003 56491
rect 44281 56457 44315 56491
rect 50169 56457 50203 56491
rect 51457 56457 51491 56491
rect 52837 56457 52871 56491
rect 53849 56457 53883 56491
rect 26341 56389 26375 56423
rect 28089 56389 28123 56423
rect 28273 56389 28307 56423
rect 33057 56389 33091 56423
rect 39865 56389 39899 56423
rect 43913 56389 43947 56423
rect 22661 56321 22695 56355
rect 23397 56321 23431 56355
rect 24041 56321 24075 56355
rect 24225 56321 24259 56355
rect 25421 56321 25455 56355
rect 26065 56321 26099 56355
rect 27169 56321 27203 56355
rect 29653 56321 29687 56355
rect 31125 56321 31159 56355
rect 32229 56321 32263 56355
rect 33241 56321 33275 56355
rect 34161 56321 34195 56355
rect 34437 56321 34471 56355
rect 35633 56321 35667 56355
rect 35817 56321 35851 56355
rect 36001 56321 36035 56355
rect 37381 56321 37415 56355
rect 39773 56321 39807 56355
rect 39957 56321 39991 56355
rect 40095 56321 40129 56355
rect 41153 56321 41187 56355
rect 42073 56321 42107 56355
rect 43269 56321 43303 56355
rect 44097 56321 44131 56355
rect 44373 56321 44407 56355
rect 45139 56321 45173 56355
rect 45293 56321 45327 56355
rect 47041 56321 47075 56355
rect 47685 56321 47719 56355
rect 48881 56321 48915 56355
rect 49525 56321 49559 56355
rect 24409 56253 24443 56287
rect 25605 56253 25639 56287
rect 27353 56253 27387 56287
rect 29837 56253 29871 56287
rect 30941 56253 30975 56287
rect 31033 56253 31067 56287
rect 31217 56253 31251 56287
rect 32505 56253 32539 56287
rect 33517 56253 33551 56287
rect 34345 56253 34379 56287
rect 34989 56253 35023 56287
rect 37473 56253 37507 56287
rect 38025 56253 38059 56287
rect 38485 56253 38519 56287
rect 40233 56253 40267 56287
rect 41429 56253 41463 56287
rect 42349 56253 42383 56287
rect 43361 56253 43395 56287
rect 46397 56253 46431 56287
rect 38117 56185 38151 56219
rect 41889 56185 41923 56219
rect 42901 56185 42935 56219
rect 45753 56185 45787 56219
rect 25237 56117 25271 56151
rect 26985 56117 27019 56151
rect 29469 56117 29503 56151
rect 30757 56117 30791 56151
rect 32413 56117 32447 56151
rect 33425 56117 33459 56151
rect 38945 56117 38979 56151
rect 41337 56117 41371 56151
rect 42257 56117 42291 56151
rect 45109 56117 45143 56151
rect 23949 55913 23983 55947
rect 24777 55913 24811 55947
rect 26065 55913 26099 55947
rect 27353 55913 27387 55947
rect 35081 55913 35115 55947
rect 37381 55913 37415 55947
rect 37841 55913 37875 55947
rect 41613 55913 41647 55947
rect 44281 55913 44315 55947
rect 45017 55913 45051 55947
rect 45661 55913 45695 55947
rect 47593 55913 47627 55947
rect 48329 55913 48363 55947
rect 25421 55845 25455 55879
rect 28641 55845 28675 55879
rect 31033 55845 31067 55879
rect 33057 55845 33091 55879
rect 39773 55845 39807 55879
rect 43637 55845 43671 55879
rect 27813 55777 27847 55811
rect 29009 55777 29043 55811
rect 31677 55777 31711 55811
rect 35449 55777 35483 55811
rect 36369 55777 36403 55811
rect 42257 55777 42291 55811
rect 43545 55777 43579 55811
rect 24593 55709 24627 55743
rect 25881 55709 25915 55743
rect 27077 55709 27111 55743
rect 27169 55709 27203 55743
rect 28825 55709 28859 55743
rect 28917 55709 28951 55743
rect 29101 55709 29135 55743
rect 30297 55709 30331 55743
rect 30481 55709 30515 55743
rect 31218 55719 31252 55753
rect 31401 55709 31435 55743
rect 32321 55709 32355 55743
rect 32597 55709 32631 55743
rect 33260 55709 33294 55743
rect 33517 55709 33551 55743
rect 34344 55709 34378 55743
rect 34437 55709 34471 55743
rect 35279 55709 35313 55743
rect 36553 55709 36587 55743
rect 36829 55709 36863 55743
rect 38025 55709 38059 55743
rect 38117 55709 38151 55743
rect 38301 55709 38335 55743
rect 38393 55709 38427 55743
rect 40601 55709 40635 55743
rect 40877 55709 40911 55743
rect 41797 55709 41831 55743
rect 43453 55709 43487 55743
rect 43729 55709 43763 55743
rect 44557 55709 44591 55743
rect 27353 55641 27387 55675
rect 27997 55641 28031 55675
rect 28181 55641 28215 55675
rect 30113 55641 30147 55675
rect 31309 55641 31343 55675
rect 31539 55641 31573 55675
rect 32505 55641 32539 55675
rect 38945 55641 38979 55675
rect 39129 55641 39163 55675
rect 39313 55641 39347 55675
rect 40785 55641 40819 55675
rect 43269 55641 43303 55675
rect 44281 55641 44315 55675
rect 44465 55641 44499 55675
rect 23489 55573 23523 55607
rect 32137 55573 32171 55607
rect 33425 55573 33459 55607
rect 34069 55573 34103 55607
rect 36737 55573 36771 55607
rect 40417 55573 40451 55607
rect 41337 55573 41371 55607
rect 46949 55573 46983 55607
rect 25329 55369 25363 55403
rect 25973 55369 26007 55403
rect 26801 55369 26835 55403
rect 27445 55369 27479 55403
rect 28549 55369 28583 55403
rect 30481 55369 30515 55403
rect 31309 55369 31343 55403
rect 35547 55369 35581 55403
rect 35633 55369 35667 55403
rect 37295 55369 37329 55403
rect 37933 55369 37967 55403
rect 38301 55369 38335 55403
rect 39957 55369 39991 55403
rect 41137 55369 41171 55403
rect 41797 55369 41831 55403
rect 46213 55369 46247 55403
rect 28089 55301 28123 55335
rect 34989 55301 35023 55335
rect 35449 55301 35483 55335
rect 37197 55301 37231 55335
rect 41337 55301 41371 55335
rect 25513 55233 25547 55267
rect 26157 55233 26191 55267
rect 26617 55233 26651 55267
rect 27261 55233 27295 55267
rect 29469 55233 29503 55267
rect 29561 55233 29595 55267
rect 29745 55233 29779 55267
rect 29837 55233 29871 55267
rect 30297 55233 30331 55267
rect 30941 55233 30975 55267
rect 31125 55233 31159 55267
rect 31953 55233 31987 55267
rect 33517 55233 33551 55267
rect 34529 55233 34563 55267
rect 34805 55233 34839 55267
rect 35725 55233 35759 55267
rect 37381 55233 37415 55267
rect 37473 55233 37507 55267
rect 38117 55233 38151 55267
rect 38393 55233 38427 55267
rect 39037 55233 39071 55267
rect 40417 55233 40451 55267
rect 42073 55233 42107 55267
rect 43269 55233 43303 55267
rect 44097 55233 44131 55267
rect 45109 55233 45143 55267
rect 45569 55233 45603 55267
rect 29285 55165 29319 55199
rect 36185 55165 36219 55199
rect 38945 55165 38979 55199
rect 41981 55165 42015 55199
rect 42441 55165 42475 55199
rect 43361 55165 43395 55199
rect 43913 55165 43947 55199
rect 44373 55165 44407 55199
rect 28457 55097 28491 55131
rect 34621 55097 34655 55131
rect 34713 55097 34747 55131
rect 42901 55097 42935 55131
rect 44281 55097 44315 55131
rect 24041 55029 24075 55063
rect 24593 55029 24627 55063
rect 32045 55029 32079 55063
rect 32413 55029 32447 55063
rect 33057 55029 33091 55063
rect 33425 55029 33459 55063
rect 39405 55029 39439 55063
rect 40325 55029 40359 55063
rect 40969 55029 41003 55063
rect 41153 55029 41187 55063
rect 44925 55029 44959 55063
rect 25421 54825 25455 54859
rect 27721 54825 27755 54859
rect 28365 54825 28399 54859
rect 31033 54825 31067 54859
rect 33149 54825 33183 54859
rect 35909 54825 35943 54859
rect 36553 54825 36587 54859
rect 37197 54825 37231 54859
rect 38025 54825 38059 54859
rect 38945 54825 38979 54859
rect 40141 54825 40175 54859
rect 42257 54825 42291 54859
rect 42901 54825 42935 54859
rect 43545 54825 43579 54859
rect 29377 54757 29411 54791
rect 32689 54757 32723 54791
rect 29101 54689 29135 54723
rect 31493 54689 31527 54723
rect 32413 54689 32447 54723
rect 33885 54689 33919 54723
rect 38393 54689 38427 54723
rect 40877 54689 40911 54723
rect 28181 54621 28215 54655
rect 28365 54621 28399 54655
rect 29009 54621 29043 54655
rect 30297 54621 30331 54655
rect 30481 54621 30515 54655
rect 31401 54621 31435 54655
rect 32321 54621 32355 54655
rect 33977 54621 34011 54655
rect 34345 54621 34379 54655
rect 35173 54621 35207 54655
rect 35265 54621 35299 54655
rect 35357 54621 35391 54655
rect 36093 54621 36127 54655
rect 38209 54621 38243 54655
rect 39129 54621 39163 54655
rect 39221 54621 39255 54655
rect 39957 54621 39991 54655
rect 40969 54621 41003 54655
rect 41797 54621 41831 54655
rect 41889 54621 41923 54655
rect 42073 54621 42107 54655
rect 39773 54553 39807 54587
rect 24593 54485 24627 54519
rect 26433 54485 26467 54519
rect 30113 54485 30147 54519
rect 33701 54485 33735 54519
rect 34989 54485 35023 54519
rect 41337 54485 41371 54519
rect 25881 54281 25915 54315
rect 26433 54281 26467 54315
rect 27353 54281 27387 54315
rect 29561 54281 29595 54315
rect 30113 54281 30147 54315
rect 31033 54281 31067 54315
rect 32413 54281 32447 54315
rect 33517 54281 33551 54315
rect 35541 54281 35575 54315
rect 38209 54281 38243 54315
rect 39589 54281 39623 54315
rect 41153 54281 41187 54315
rect 41797 54281 41831 54315
rect 42809 54281 42843 54315
rect 29377 54213 29411 54247
rect 30481 54213 30515 54247
rect 31217 54213 31251 54247
rect 37657 54213 37691 54247
rect 38393 54213 38427 54247
rect 38577 54213 38611 54247
rect 39773 54213 39807 54247
rect 27905 54145 27939 54179
rect 28365 54145 28399 54179
rect 29653 54145 29687 54179
rect 30297 54145 30331 54179
rect 30941 54145 30975 54179
rect 32229 54145 32263 54179
rect 32505 54145 32539 54179
rect 33885 54145 33919 54179
rect 34713 54145 34747 54179
rect 34989 54145 35023 54179
rect 35633 54145 35667 54179
rect 36093 54145 36127 54179
rect 37013 54145 37047 54179
rect 39497 54145 39531 54179
rect 40969 54145 41003 54179
rect 41985 54145 42019 54179
rect 42083 54151 42117 54185
rect 42201 54145 42235 54179
rect 32045 54077 32079 54111
rect 33977 54077 34011 54111
rect 34529 54077 34563 54111
rect 34897 54077 34931 54111
rect 29377 54009 29411 54043
rect 31217 54009 31251 54043
rect 39773 54009 39807 54043
rect 28549 53941 28583 53975
rect 40233 53941 40267 53975
rect 28181 53737 28215 53771
rect 29285 53737 29319 53771
rect 30021 53737 30055 53771
rect 32689 53737 32723 53771
rect 33609 53737 33643 53771
rect 33793 53737 33827 53771
rect 35725 53737 35759 53771
rect 36829 53737 36863 53771
rect 37841 53737 37875 53771
rect 38945 53737 38979 53771
rect 39681 53737 39715 53771
rect 40233 53737 40267 53771
rect 40785 53737 40819 53771
rect 41429 53737 41463 53771
rect 36369 53669 36403 53703
rect 28825 53601 28859 53635
rect 29285 53533 29319 53567
rect 29469 53533 29503 53567
rect 32873 53533 32907 53567
rect 33057 53533 33091 53567
rect 33149 53533 33183 53567
rect 35173 53533 35207 53567
rect 39773 53533 39807 53567
rect 33772 53465 33806 53499
rect 33977 53465 34011 53499
rect 31401 53397 31435 53431
rect 31953 53397 31987 53431
rect 30297 53193 30331 53227
rect 33701 53193 33735 53227
rect 39037 53193 39071 53227
rect 39957 53193 39991 53227
rect 40969 53193 41003 53227
rect 33149 53125 33183 53159
rect 35909 53125 35943 53159
rect 38577 53125 38611 53159
rect 29561 53057 29595 53091
rect 36093 53057 36127 53091
rect 34529 52989 34563 53023
rect 29377 52649 29411 52683
rect 35081 52649 35115 52683
rect 36093 52649 36127 52683
rect 26433 8041 26467 8075
rect 25973 7429 26007 7463
rect 29653 7361 29687 7395
rect 25789 7293 25823 7327
rect 26801 7293 26835 7327
rect 28089 7157 28123 7191
rect 29745 7157 29779 7191
rect 30389 7157 30423 7191
rect 27997 6817 28031 6851
rect 28641 6817 28675 6851
rect 25973 6749 26007 6783
rect 27353 6749 27387 6783
rect 30297 6749 30331 6783
rect 31033 6749 31067 6783
rect 32137 6749 32171 6783
rect 26525 6681 26559 6715
rect 28181 6681 28215 6715
rect 25881 6613 25915 6647
rect 27445 6613 27479 6647
rect 32229 6613 32263 6647
rect 26157 6341 26191 6375
rect 26893 6341 26927 6375
rect 29745 6341 29779 6375
rect 35633 6341 35667 6375
rect 26065 6273 26099 6307
rect 29561 6273 29595 6307
rect 31861 6273 31895 6307
rect 26709 6205 26743 6239
rect 27905 6205 27939 6239
rect 30205 6205 30239 6239
rect 34437 6205 34471 6239
rect 35817 6205 35851 6239
rect 24041 6069 24075 6103
rect 25421 6069 25455 6103
rect 31953 6069 31987 6103
rect 33057 6069 33091 6103
rect 24685 5729 24719 5763
rect 24869 5729 24903 5763
rect 26157 5729 26191 5763
rect 28089 5729 28123 5763
rect 30297 5729 30331 5763
rect 31033 5729 31067 5763
rect 31217 5729 31251 5763
rect 31677 5729 31711 5763
rect 23213 5661 23247 5695
rect 24225 5661 24259 5695
rect 27537 5661 27571 5695
rect 30021 5661 30055 5695
rect 33333 5661 33367 5695
rect 34161 5661 34195 5695
rect 35173 5661 35207 5695
rect 27721 5593 27755 5627
rect 24133 5525 24167 5559
rect 34069 5525 34103 5559
rect 35081 5525 35115 5559
rect 25237 5321 25271 5355
rect 22937 5253 22971 5287
rect 26893 5253 26927 5287
rect 34805 5253 34839 5287
rect 25145 5185 25179 5219
rect 25789 5185 25823 5219
rect 26709 5185 26743 5219
rect 22753 5117 22787 5151
rect 24593 5117 24627 5151
rect 25973 5117 26007 5151
rect 28365 5117 28399 5151
rect 29653 5117 29687 5151
rect 30113 5117 30147 5151
rect 30297 5117 30331 5151
rect 30573 5117 30607 5151
rect 33333 5117 33367 5151
rect 34989 5117 35023 5151
rect 35449 5117 35483 5151
rect 22293 4981 22327 5015
rect 32413 4981 32447 5015
rect 36093 4981 36127 5015
rect 22569 4777 22603 4811
rect 27537 4777 27571 4811
rect 21925 4709 21959 4743
rect 37933 4709 37967 4743
rect 30021 4641 30055 4675
rect 31309 4641 31343 4675
rect 32045 4641 32079 4675
rect 32229 4641 32263 4675
rect 32781 4641 32815 4675
rect 19349 4573 19383 4607
rect 20453 4573 20487 4607
rect 21281 4573 21315 4607
rect 23397 4573 23431 4607
rect 24225 4573 24259 4607
rect 24685 4573 24719 4607
rect 28181 4573 28215 4607
rect 28641 4573 28675 4607
rect 31033 4573 31067 4607
rect 36829 4573 36863 4607
rect 37289 4573 37323 4607
rect 38945 4573 38979 4607
rect 23489 4505 23523 4539
rect 24869 4505 24903 4539
rect 26525 4505 26559 4539
rect 28825 4505 28859 4539
rect 34989 4505 35023 4539
rect 36645 4505 36679 4539
rect 30113 4233 30147 4267
rect 22293 4097 22327 4131
rect 25605 4097 25639 4131
rect 26249 4097 26283 4131
rect 29377 4097 29411 4131
rect 30021 4097 30055 4131
rect 33057 4097 33091 4131
rect 35357 4097 35391 4131
rect 36185 4097 36219 4131
rect 19993 4029 20027 4063
rect 22753 4029 22787 4063
rect 22937 4029 22971 4063
rect 24593 4029 24627 4063
rect 26709 4029 26743 4063
rect 26893 4029 26927 4063
rect 28549 4029 28583 4063
rect 30665 4029 30699 4063
rect 30849 4029 30883 4063
rect 31401 4029 31435 4063
rect 33241 4029 33275 4063
rect 33517 4029 33551 4063
rect 37013 4029 37047 4063
rect 37197 4029 37231 4063
rect 37473 4029 37507 4063
rect 29469 3961 29503 3995
rect 39957 3961 39991 3995
rect 16405 3893 16439 3927
rect 17693 3893 17727 3927
rect 18521 3893 18555 3927
rect 19349 3893 19383 3927
rect 20637 3893 20671 3927
rect 21649 3893 21683 3927
rect 35449 3893 35483 3927
rect 39313 3893 39347 3927
rect 40969 3893 41003 3927
rect 23397 3689 23431 3723
rect 27445 3689 27479 3723
rect 27997 3689 28031 3723
rect 31033 3689 31067 3723
rect 37381 3689 37415 3723
rect 37933 3689 37967 3723
rect 39589 3689 39623 3723
rect 19625 3621 19659 3655
rect 38945 3621 38979 3655
rect 40877 3621 40911 3655
rect 42901 3621 42935 3655
rect 44189 3621 44223 3655
rect 46121 3621 46155 3655
rect 18613 3553 18647 3587
rect 22017 3553 22051 3587
rect 26065 3553 26099 3587
rect 28641 3553 28675 3587
rect 32505 3553 32539 3587
rect 35449 3553 35483 3587
rect 40233 3553 40267 3587
rect 41521 3553 41555 3587
rect 44833 3553 44867 3587
rect 9413 3485 9447 3519
rect 10333 3485 10367 3519
rect 11989 3485 12023 3519
rect 12817 3485 12851 3519
rect 13645 3485 13679 3519
rect 14473 3485 14507 3519
rect 15209 3485 15243 3519
rect 15853 3485 15887 3519
rect 16681 3485 16715 3519
rect 17325 3485 17359 3519
rect 17969 3485 18003 3519
rect 20269 3485 20303 3519
rect 22569 3485 22603 3519
rect 24225 3485 24259 3519
rect 26525 3485 26559 3519
rect 27537 3485 27571 3519
rect 33701 3485 33735 3519
rect 34345 3485 34379 3519
rect 34989 3485 35023 3519
rect 37473 3485 37507 3519
rect 42165 3485 42199 3519
rect 43545 3485 43579 3519
rect 45477 3485 45511 3519
rect 46857 3485 46891 3519
rect 47501 3485 47535 3519
rect 48145 3485 48179 3519
rect 49157 3485 49191 3519
rect 49801 3485 49835 3519
rect 51089 3485 51123 3519
rect 51733 3485 51767 3519
rect 22385 3417 22419 3451
rect 26341 3417 26375 3451
rect 28825 3417 28859 3451
rect 30481 3417 30515 3451
rect 33517 3417 33551 3451
rect 34253 3417 34287 3451
rect 35173 3417 35207 3451
rect 21557 3145 21591 3179
rect 29469 3145 29503 3179
rect 37197 3077 37231 3111
rect 18705 3009 18739 3043
rect 21649 3009 21683 3043
rect 22293 3009 22327 3043
rect 24593 3009 24627 3043
rect 25605 3009 25639 3043
rect 29561 3009 29595 3043
rect 35357 3009 35391 3043
rect 37013 3009 37047 3043
rect 40969 3009 41003 3043
rect 42901 3009 42935 3043
rect 15393 2941 15427 2975
rect 17417 2941 17451 2975
rect 19349 2941 19383 2975
rect 24133 2941 24167 2975
rect 24409 2941 24443 2975
rect 26249 2941 26283 2975
rect 26709 2941 26743 2975
rect 26893 2941 26927 2975
rect 28549 2941 28583 2975
rect 30113 2941 30147 2975
rect 30297 2941 30331 2975
rect 31217 2941 31251 2975
rect 33057 2941 33091 2975
rect 34713 2941 34747 2975
rect 34897 2941 34931 2975
rect 36185 2941 36219 2975
rect 37657 2941 37691 2975
rect 41613 2941 41647 2975
rect 43545 2941 43579 2975
rect 45569 2941 45603 2975
rect 47501 2941 47535 2975
rect 50813 2941 50847 2975
rect 52837 2941 52871 2975
rect 18061 2873 18095 2907
rect 19993 2873 20027 2907
rect 20637 2873 20671 2907
rect 39957 2873 39991 2907
rect 42257 2873 42291 2907
rect 44189 2873 44223 2907
rect 46213 2873 46247 2907
rect 48145 2873 48179 2907
rect 49525 2873 49559 2907
rect 51457 2873 51491 2907
rect 7481 2805 7515 2839
rect 8125 2805 8159 2839
rect 8769 2805 8803 2839
rect 9505 2805 9539 2839
rect 10149 2805 10183 2839
rect 10793 2805 10827 2839
rect 11437 2805 11471 2839
rect 12081 2805 12115 2839
rect 12725 2805 12759 2839
rect 13461 2805 13495 2839
rect 14105 2805 14139 2839
rect 14749 2805 14783 2839
rect 16037 2805 16071 2839
rect 16681 2805 16715 2839
rect 39313 2805 39347 2839
rect 44925 2805 44959 2839
rect 46857 2805 46891 2839
rect 48881 2805 48915 2839
rect 50169 2805 50203 2839
rect 52101 2805 52135 2839
rect 23305 2601 23339 2635
rect 23949 2601 23983 2635
rect 25237 2601 25271 2635
rect 27169 2601 27203 2635
rect 27813 2601 27847 2635
rect 29101 2601 29135 2635
rect 29653 2601 29687 2635
rect 30389 2601 30423 2635
rect 31125 2601 31159 2635
rect 32505 2601 32539 2635
rect 34345 2601 34379 2635
rect 34989 2601 35023 2635
rect 36369 2601 36403 2635
rect 38209 2601 38243 2635
rect 38761 2601 38795 2635
rect 40049 2601 40083 2635
rect 7941 2533 7975 2567
rect 11805 2533 11839 2567
rect 16313 2533 16347 2567
rect 21465 2533 21499 2567
rect 33149 2533 33183 2567
rect 36921 2533 36955 2567
rect 42625 2533 42659 2567
rect 45845 2533 45879 2567
rect 48421 2533 48455 2567
rect 53573 2533 53607 2567
rect 9873 2465 9907 2499
rect 13737 2465 13771 2499
rect 15669 2465 15703 2499
rect 17601 2465 17635 2499
rect 22109 2465 22143 2499
rect 41981 2465 42015 2499
rect 44557 2465 44591 2499
rect 46489 2465 46523 2499
rect 49709 2465 49743 2499
rect 51641 2465 51675 2499
rect 54217 2465 54251 2499
rect 8585 2397 8619 2431
rect 10517 2397 10551 2431
rect 12449 2397 12483 2431
rect 14381 2397 14415 2431
rect 18245 2397 18279 2431
rect 19533 2397 19567 2431
rect 20177 2397 20211 2431
rect 23397 2397 23431 2431
rect 24041 2397 24075 2431
rect 25329 2397 25363 2431
rect 25789 2397 25823 2431
rect 27261 2397 27295 2431
rect 27905 2397 27939 2431
rect 29193 2397 29227 2431
rect 31217 2397 31251 2431
rect 34437 2397 34471 2431
rect 34897 2397 34931 2431
rect 36829 2397 36863 2431
rect 38117 2397 38151 2431
rect 40693 2397 40727 2431
rect 43913 2397 43947 2431
rect 47777 2397 47811 2431
rect 50353 2397 50387 2431
rect 52285 2397 52319 2431
rect 25881 2329 25915 2363
<< metal1 >>
rect 15194 57876 15200 57928
rect 15252 57916 15258 57928
rect 25682 57916 25688 57928
rect 15252 57888 25688 57916
rect 15252 57876 15258 57888
rect 25682 57876 25688 57888
rect 25740 57876 25746 57928
rect 27614 57876 27620 57928
rect 27672 57916 27678 57928
rect 35986 57916 35992 57928
rect 27672 57888 35992 57916
rect 27672 57876 27678 57888
rect 35986 57876 35992 57888
rect 36044 57876 36050 57928
rect 22002 57808 22008 57860
rect 22060 57848 22066 57860
rect 24670 57848 24676 57860
rect 22060 57820 24676 57848
rect 22060 57808 22066 57820
rect 24670 57808 24676 57820
rect 24728 57808 24734 57860
rect 24762 57808 24768 57860
rect 24820 57848 24826 57860
rect 40034 57848 40040 57860
rect 24820 57820 40040 57848
rect 24820 57808 24826 57820
rect 40034 57808 40040 57820
rect 40092 57808 40098 57860
rect 40126 57808 40132 57860
rect 40184 57848 40190 57860
rect 40184 57820 40540 57848
rect 40184 57808 40190 57820
rect 20990 57740 20996 57792
rect 21048 57780 21054 57792
rect 25038 57780 25044 57792
rect 21048 57752 25044 57780
rect 21048 57740 21054 57752
rect 25038 57740 25044 57752
rect 25096 57740 25102 57792
rect 27982 57740 27988 57792
rect 28040 57780 28046 57792
rect 35526 57780 35532 57792
rect 28040 57752 35532 57780
rect 28040 57740 28046 57752
rect 35526 57740 35532 57752
rect 35584 57740 35590 57792
rect 35710 57740 35716 57792
rect 35768 57780 35774 57792
rect 40402 57780 40408 57792
rect 35768 57752 40408 57780
rect 35768 57740 35774 57752
rect 40402 57740 40408 57752
rect 40460 57740 40466 57792
rect 40512 57780 40540 57820
rect 42334 57808 42340 57860
rect 42392 57848 42398 57860
rect 44726 57848 44732 57860
rect 42392 57820 44732 57848
rect 42392 57808 42398 57820
rect 44726 57808 44732 57820
rect 44784 57808 44790 57860
rect 49142 57780 49148 57792
rect 40512 57752 49148 57780
rect 49142 57740 49148 57752
rect 49200 57740 49206 57792
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 5074 57536 5080 57588
rect 5132 57576 5138 57588
rect 5353 57579 5411 57585
rect 5353 57576 5365 57579
rect 5132 57548 5365 57576
rect 5132 57536 5138 57548
rect 5353 57545 5365 57548
rect 5399 57545 5411 57579
rect 5353 57539 5411 57545
rect 11054 57536 11060 57588
rect 11112 57576 11118 57588
rect 11149 57579 11207 57585
rect 11149 57576 11161 57579
rect 11112 57548 11161 57576
rect 11112 57536 11118 57548
rect 11149 57545 11161 57548
rect 11195 57545 11207 57579
rect 11149 57539 11207 57545
rect 11974 57536 11980 57588
rect 12032 57576 12038 57588
rect 12161 57579 12219 57585
rect 12161 57576 12173 57579
rect 12032 57548 12173 57576
rect 12032 57536 12038 57548
rect 12161 57545 12173 57548
rect 12207 57545 12219 57579
rect 12161 57539 12219 57545
rect 13354 57536 13360 57588
rect 13412 57576 13418 57588
rect 13541 57579 13599 57585
rect 13541 57576 13553 57579
rect 13412 57548 13553 57576
rect 13412 57536 13418 57548
rect 13541 57545 13553 57548
rect 13587 57545 13599 57579
rect 13541 57539 13599 57545
rect 14734 57536 14740 57588
rect 14792 57576 14798 57588
rect 15013 57579 15071 57585
rect 15013 57576 15025 57579
rect 14792 57548 15025 57576
rect 14792 57536 14798 57548
rect 15013 57545 15025 57548
rect 15059 57545 15071 57579
rect 15013 57539 15071 57545
rect 16114 57536 16120 57588
rect 16172 57576 16178 57588
rect 16945 57579 17003 57585
rect 16945 57576 16957 57579
rect 16172 57548 16957 57576
rect 16172 57536 16178 57548
rect 16945 57545 16957 57548
rect 16991 57545 17003 57579
rect 16945 57539 17003 57545
rect 17494 57536 17500 57588
rect 17552 57576 17558 57588
rect 17681 57579 17739 57585
rect 17681 57576 17693 57579
rect 17552 57548 17693 57576
rect 17552 57536 17558 57548
rect 17681 57545 17693 57548
rect 17727 57545 17739 57579
rect 17681 57539 17739 57545
rect 18874 57536 18880 57588
rect 18932 57576 18938 57588
rect 19061 57579 19119 57585
rect 19061 57576 19073 57579
rect 18932 57548 19073 57576
rect 18932 57536 18938 57548
rect 19061 57545 19073 57548
rect 19107 57545 19119 57579
rect 19061 57539 19119 57545
rect 20254 57536 20260 57588
rect 20312 57576 20318 57588
rect 20809 57579 20867 57585
rect 20809 57576 20821 57579
rect 20312 57548 20821 57576
rect 20312 57536 20318 57548
rect 20809 57545 20821 57548
rect 20855 57545 20867 57579
rect 20809 57539 20867 57545
rect 21634 57536 21640 57588
rect 21692 57576 21698 57588
rect 21821 57579 21879 57585
rect 21821 57576 21833 57579
rect 21692 57548 21833 57576
rect 21692 57536 21698 57548
rect 21821 57545 21833 57548
rect 21867 57545 21879 57579
rect 21821 57539 21879 57545
rect 23014 57536 23020 57588
rect 23072 57576 23078 57588
rect 23109 57579 23167 57585
rect 23109 57576 23121 57579
rect 23072 57548 23121 57576
rect 23072 57536 23078 57548
rect 23109 57545 23121 57548
rect 23155 57545 23167 57579
rect 23109 57539 23167 57545
rect 23937 57579 23995 57585
rect 23937 57545 23949 57579
rect 23983 57576 23995 57579
rect 24394 57576 24400 57588
rect 23983 57548 24400 57576
rect 23983 57545 23995 57548
rect 23937 57539 23995 57545
rect 24394 57536 24400 57548
rect 24452 57536 24458 57588
rect 24670 57536 24676 57588
rect 24728 57576 24734 57588
rect 25958 57576 25964 57588
rect 24728 57548 25964 57576
rect 24728 57536 24734 57548
rect 25958 57536 25964 57548
rect 26016 57576 26022 57588
rect 27062 57576 27068 57588
rect 26016 57548 27068 57576
rect 26016 57536 26022 57548
rect 27062 57536 27068 57548
rect 27120 57536 27126 57588
rect 31294 57536 31300 57588
rect 31352 57576 31358 57588
rect 34238 57576 34244 57588
rect 31352 57548 34244 57576
rect 31352 57536 31358 57548
rect 34238 57536 34244 57548
rect 34296 57536 34302 57588
rect 40034 57576 40040 57588
rect 39995 57548 40040 57576
rect 40034 57536 40040 57548
rect 40092 57536 40098 57588
rect 41969 57579 42027 57585
rect 41969 57576 41981 57579
rect 40144 57548 41981 57576
rect 3694 57468 3700 57520
rect 3752 57508 3758 57520
rect 3881 57511 3939 57517
rect 3881 57508 3893 57511
rect 3752 57480 3893 57508
rect 3752 57468 3758 57480
rect 3881 57477 3893 57480
rect 3927 57477 3939 57511
rect 23198 57508 23204 57520
rect 3881 57471 3939 57477
rect 13740 57480 23204 57508
rect 4525 57443 4583 57449
rect 4525 57409 4537 57443
rect 4571 57440 4583 57443
rect 4614 57440 4620 57452
rect 4571 57412 4620 57440
rect 4571 57409 4583 57412
rect 4525 57403 4583 57409
rect 4614 57400 4620 57412
rect 4672 57400 4678 57452
rect 5537 57443 5595 57449
rect 5537 57409 5549 57443
rect 5583 57409 5595 57443
rect 6454 57440 6460 57452
rect 6415 57412 6460 57440
rect 5537 57403 5595 57409
rect 5552 57372 5580 57403
rect 6454 57400 6460 57412
rect 6512 57400 6518 57452
rect 7745 57443 7803 57449
rect 7745 57409 7757 57443
rect 7791 57440 7803 57443
rect 7834 57440 7840 57452
rect 7791 57412 7840 57440
rect 7791 57409 7803 57412
rect 7745 57403 7803 57409
rect 7834 57400 7840 57412
rect 7892 57400 7898 57452
rect 8573 57443 8631 57449
rect 8573 57409 8585 57443
rect 8619 57440 8631 57443
rect 8754 57440 8760 57452
rect 8619 57412 8760 57440
rect 8619 57409 8631 57412
rect 8573 57403 8631 57409
rect 8754 57400 8760 57412
rect 8812 57400 8818 57452
rect 9214 57400 9220 57452
rect 9272 57440 9278 57452
rect 9309 57443 9367 57449
rect 9309 57440 9321 57443
rect 9272 57412 9321 57440
rect 9272 57400 9278 57412
rect 9309 57409 9321 57412
rect 9355 57409 9367 57443
rect 9309 57403 9367 57409
rect 10134 57400 10140 57452
rect 10192 57440 10198 57452
rect 10229 57443 10287 57449
rect 10229 57440 10241 57443
rect 10192 57412 10241 57440
rect 10192 57400 10198 57412
rect 10229 57409 10241 57412
rect 10275 57409 10287 57443
rect 11330 57440 11336 57452
rect 11291 57412 11336 57440
rect 10229 57403 10287 57409
rect 11330 57400 11336 57412
rect 11388 57400 11394 57452
rect 12342 57440 12348 57452
rect 12303 57412 12348 57440
rect 12342 57400 12348 57412
rect 12400 57400 12406 57452
rect 13740 57449 13768 57480
rect 23198 57468 23204 57480
rect 23256 57468 23262 57520
rect 33686 57508 33692 57520
rect 23308 57480 29684 57508
rect 13725 57443 13783 57449
rect 13725 57409 13737 57443
rect 13771 57409 13783 57443
rect 13725 57403 13783 57409
rect 14185 57443 14243 57449
rect 14185 57409 14197 57443
rect 14231 57440 14243 57443
rect 14274 57440 14280 57452
rect 14231 57412 14280 57440
rect 14231 57409 14243 57412
rect 14185 57403 14243 57409
rect 14274 57400 14280 57412
rect 14332 57400 14338 57452
rect 15194 57440 15200 57452
rect 15155 57412 15200 57440
rect 15194 57400 15200 57412
rect 15252 57400 15258 57452
rect 15654 57400 15660 57452
rect 15712 57440 15718 57452
rect 15749 57443 15807 57449
rect 15749 57440 15761 57443
rect 15712 57412 15761 57440
rect 15712 57400 15718 57412
rect 15749 57409 15761 57412
rect 15795 57409 15807 57443
rect 15749 57403 15807 57409
rect 17129 57443 17187 57449
rect 17129 57409 17141 57443
rect 17175 57409 17187 57443
rect 17129 57403 17187 57409
rect 17865 57443 17923 57449
rect 17865 57409 17877 57443
rect 17911 57409 17923 57443
rect 19242 57440 19248 57452
rect 19203 57412 19248 57440
rect 17865 57403 17923 57409
rect 7282 57372 7288 57384
rect 5552 57344 7288 57372
rect 7282 57332 7288 57344
rect 7340 57332 7346 57384
rect 4065 57307 4123 57313
rect 4065 57273 4077 57307
rect 4111 57304 4123 57307
rect 16942 57304 16948 57316
rect 4111 57276 16948 57304
rect 4111 57273 4123 57276
rect 4065 57267 4123 57273
rect 16942 57264 16948 57276
rect 17000 57264 17006 57316
rect 7282 57236 7288 57248
rect 7243 57208 7288 57236
rect 7282 57196 7288 57208
rect 7340 57196 7346 57248
rect 17144 57236 17172 57403
rect 17880 57372 17908 57403
rect 19242 57400 19248 57412
rect 19300 57400 19306 57452
rect 19889 57443 19947 57449
rect 19889 57409 19901 57443
rect 19935 57440 19947 57443
rect 19978 57440 19984 57452
rect 19935 57412 19984 57440
rect 19935 57409 19947 57412
rect 19889 57403 19947 57409
rect 19978 57400 19984 57412
rect 20036 57400 20042 57452
rect 20990 57440 20996 57452
rect 20951 57412 20996 57440
rect 20990 57400 20996 57412
rect 21048 57400 21054 57452
rect 22002 57440 22008 57452
rect 21963 57412 22008 57440
rect 22002 57400 22008 57412
rect 22060 57400 22066 57452
rect 23308 57449 23336 57480
rect 23293 57443 23351 57449
rect 23293 57409 23305 57443
rect 23339 57409 23351 57443
rect 23750 57440 23756 57452
rect 23711 57412 23756 57440
rect 23293 57403 23351 57409
rect 23750 57400 23756 57412
rect 23808 57400 23814 57452
rect 24762 57440 24768 57452
rect 24723 57412 24768 57440
rect 24762 57400 24768 57412
rect 24820 57400 24826 57452
rect 25590 57440 25596 57452
rect 25551 57412 25596 57440
rect 25590 57400 25596 57412
rect 25648 57400 25654 57452
rect 26418 57400 26424 57452
rect 26476 57440 26482 57452
rect 26881 57443 26939 57449
rect 26881 57440 26893 57443
rect 26476 57412 26893 57440
rect 26476 57400 26482 57412
rect 26881 57409 26893 57412
rect 26927 57409 26939 57443
rect 26881 57403 26939 57409
rect 27157 57443 27215 57449
rect 27157 57409 27169 57443
rect 27203 57440 27215 57443
rect 27614 57440 27620 57452
rect 27203 57412 27620 57440
rect 27203 57409 27215 57412
rect 27157 57403 27215 57409
rect 27614 57400 27620 57412
rect 27672 57400 27678 57452
rect 27890 57440 27896 57452
rect 27851 57412 27896 57440
rect 27890 57400 27896 57412
rect 27948 57400 27954 57452
rect 29089 57443 29147 57449
rect 29089 57409 29101 57443
rect 29135 57440 29147 57443
rect 29178 57440 29184 57452
rect 29135 57412 29184 57440
rect 29135 57409 29147 57412
rect 29089 57403 29147 57409
rect 29178 57400 29184 57412
rect 29236 57400 29242 57452
rect 29270 57400 29276 57452
rect 29328 57440 29334 57452
rect 29549 57443 29607 57449
rect 29328 57412 29373 57440
rect 29328 57400 29334 57412
rect 29549 57409 29561 57443
rect 29595 57440 29607 57443
rect 29656 57440 29684 57480
rect 30300 57480 33692 57508
rect 30300 57440 30328 57480
rect 33686 57468 33692 57480
rect 33744 57468 33750 57520
rect 34514 57468 34520 57520
rect 34572 57508 34578 57520
rect 34701 57511 34759 57517
rect 34701 57508 34713 57511
rect 34572 57480 34713 57508
rect 34572 57468 34578 57480
rect 34701 57477 34713 57480
rect 34747 57508 34759 57511
rect 40144 57508 40172 57548
rect 41969 57545 41981 57548
rect 42015 57545 42027 57579
rect 41969 57539 42027 57545
rect 43346 57536 43352 57588
rect 43404 57576 43410 57588
rect 47995 57579 48053 57585
rect 47995 57576 48007 57579
rect 43404 57548 48007 57576
rect 43404 57536 43410 57548
rect 47995 57545 48007 57548
rect 48041 57545 48053 57579
rect 52641 57579 52699 57585
rect 52641 57576 52653 57579
rect 47995 57539 48053 57545
rect 51046 57548 52653 57576
rect 34747 57480 40172 57508
rect 34747 57477 34759 57480
rect 34701 57471 34759 57477
rect 40402 57468 40408 57520
rect 40460 57508 40466 57520
rect 51046 57508 51074 57548
rect 52641 57545 52653 57548
rect 52687 57545 52699 57579
rect 52641 57539 52699 57545
rect 40460 57480 51074 57508
rect 40460 57468 40466 57480
rect 52454 57468 52460 57520
rect 52512 57508 52518 57520
rect 52822 57508 52828 57520
rect 52512 57480 52828 57508
rect 52512 57468 52518 57480
rect 52822 57468 52828 57480
rect 52880 57508 52886 57520
rect 52917 57511 52975 57517
rect 52917 57508 52929 57511
rect 52880 57480 52929 57508
rect 52880 57468 52886 57480
rect 52917 57477 52929 57480
rect 52963 57477 52975 57511
rect 52917 57471 52975 57477
rect 29595 57412 30328 57440
rect 30377 57443 30435 57449
rect 29595 57409 29607 57412
rect 29549 57403 29607 57409
rect 30377 57409 30389 57443
rect 30423 57409 30435 57443
rect 31386 57440 31392 57452
rect 31347 57412 31392 57440
rect 30377 57403 30435 57409
rect 24949 57375 25007 57381
rect 17880 57344 24900 57372
rect 21358 57264 21364 57316
rect 21416 57304 21422 57316
rect 24872 57304 24900 57344
rect 24949 57341 24961 57375
rect 24995 57372 25007 57375
rect 25777 57375 25835 57381
rect 25777 57372 25789 57375
rect 24995 57344 25789 57372
rect 24995 57341 25007 57344
rect 24949 57335 25007 57341
rect 25777 57341 25789 57344
rect 25823 57372 25835 57375
rect 26142 57372 26148 57384
rect 25823 57344 26148 57372
rect 25823 57341 25835 57344
rect 25777 57335 25835 57341
rect 26142 57332 26148 57344
rect 26200 57332 26206 57384
rect 27724 57344 28396 57372
rect 27724 57304 27752 57344
rect 21416 57276 24808 57304
rect 24872 57276 27752 57304
rect 27801 57307 27859 57313
rect 21416 57264 21422 57276
rect 22462 57236 22468 57248
rect 17144 57208 22468 57236
rect 22462 57196 22468 57208
rect 22520 57196 22526 57248
rect 22646 57196 22652 57248
rect 22704 57236 22710 57248
rect 24581 57239 24639 57245
rect 24581 57236 24593 57239
rect 22704 57208 24593 57236
rect 22704 57196 22710 57208
rect 24581 57205 24593 57208
rect 24627 57205 24639 57239
rect 24780 57236 24808 57276
rect 27801 57273 27813 57307
rect 27847 57304 27859 57307
rect 28258 57304 28264 57316
rect 27847 57276 28264 57304
rect 27847 57273 27859 57276
rect 27801 57267 27859 57273
rect 28258 57264 28264 57276
rect 28316 57264 28322 57316
rect 28368 57304 28396 57344
rect 28534 57332 28540 57384
rect 28592 57372 28598 57384
rect 29365 57375 29423 57381
rect 28592 57344 29316 57372
rect 28592 57332 28598 57344
rect 28905 57307 28963 57313
rect 28905 57304 28917 57307
rect 28368 57276 28917 57304
rect 28905 57273 28917 57276
rect 28951 57273 28963 57307
rect 28905 57267 28963 57273
rect 29181 57307 29239 57313
rect 29181 57273 29193 57307
rect 29227 57273 29239 57307
rect 29288 57304 29316 57344
rect 29365 57341 29377 57375
rect 29411 57372 29423 57375
rect 30006 57372 30012 57384
rect 29411 57344 30012 57372
rect 29411 57341 29423 57344
rect 29365 57335 29423 57341
rect 30006 57332 30012 57344
rect 30064 57372 30070 57384
rect 30392 57372 30420 57403
rect 31386 57400 31392 57412
rect 31444 57400 31450 57452
rect 31754 57400 31760 57452
rect 31812 57440 31818 57452
rect 32309 57443 32367 57449
rect 32309 57440 32321 57443
rect 31812 57412 32321 57440
rect 31812 57400 31818 57412
rect 32309 57409 32321 57412
rect 32355 57440 32367 57443
rect 37461 57443 37519 57449
rect 37461 57440 37473 57443
rect 32355 57412 37473 57440
rect 32355 57409 32367 57412
rect 32309 57403 32367 57409
rect 37461 57409 37473 57412
rect 37507 57409 37519 57443
rect 37461 57403 37519 57409
rect 37550 57400 37556 57452
rect 37608 57440 37614 57452
rect 39485 57443 39543 57449
rect 39485 57440 39497 57443
rect 37608 57412 39497 57440
rect 37608 57400 37614 57412
rect 39485 57409 39497 57412
rect 39531 57440 39543 57443
rect 40126 57440 40132 57452
rect 39531 57412 40132 57440
rect 39531 57409 39543 57412
rect 39485 57403 39543 57409
rect 40126 57400 40132 57412
rect 40184 57400 40190 57452
rect 40221 57443 40279 57449
rect 40221 57409 40233 57443
rect 40267 57440 40279 57443
rect 40862 57440 40868 57452
rect 40267 57412 40868 57440
rect 40267 57409 40279 57412
rect 40221 57403 40279 57409
rect 40862 57400 40868 57412
rect 40920 57400 40926 57452
rect 41230 57440 41236 57452
rect 41191 57412 41236 57440
rect 41230 57400 41236 57412
rect 41288 57400 41294 57452
rect 41322 57400 41328 57452
rect 41380 57440 41386 57452
rect 41417 57443 41475 57449
rect 41417 57440 41429 57443
rect 41380 57412 41429 57440
rect 41380 57400 41386 57412
rect 41417 57409 41429 57412
rect 41463 57409 41475 57443
rect 41417 57403 41475 57409
rect 31662 57372 31668 57384
rect 30064 57344 30420 57372
rect 31623 57344 31668 57372
rect 30064 57332 30070 57344
rect 31662 57332 31668 57344
rect 31720 57332 31726 57384
rect 32582 57372 32588 57384
rect 32543 57344 32588 57372
rect 32582 57332 32588 57344
rect 32640 57332 32646 57384
rect 33134 57332 33140 57384
rect 33192 57372 33198 57384
rect 35802 57372 35808 57384
rect 33192 57344 35808 57372
rect 33192 57332 33198 57344
rect 35802 57332 35808 57344
rect 35860 57332 35866 57384
rect 35894 57332 35900 57384
rect 35952 57372 35958 57384
rect 36170 57372 36176 57384
rect 35952 57344 36176 57372
rect 35952 57332 35958 57344
rect 36170 57332 36176 57344
rect 36228 57332 36234 57384
rect 36449 57375 36507 57381
rect 36449 57341 36461 57375
rect 36495 57341 36507 57375
rect 36449 57335 36507 57341
rect 30561 57307 30619 57313
rect 30561 57304 30573 57307
rect 29288 57276 30573 57304
rect 29181 57267 29239 57273
rect 30561 57273 30573 57276
rect 30607 57273 30619 57307
rect 30561 57267 30619 57273
rect 25222 57236 25228 57248
rect 24780 57208 25228 57236
rect 24581 57199 24639 57205
rect 25222 57196 25228 57208
rect 25280 57196 25286 57248
rect 25409 57239 25467 57245
rect 25409 57205 25421 57239
rect 25455 57236 25467 57239
rect 25498 57236 25504 57248
rect 25455 57208 25504 57236
rect 25455 57205 25467 57208
rect 25409 57199 25467 57205
rect 25498 57196 25504 57208
rect 25556 57196 25562 57248
rect 27706 57236 27712 57248
rect 27667 57208 27712 57236
rect 27706 57196 27712 57208
rect 27764 57196 27770 57248
rect 28350 57196 28356 57248
rect 28408 57236 28414 57248
rect 29196 57236 29224 57267
rect 34422 57264 34428 57316
rect 34480 57304 34486 57316
rect 36464 57304 36492 57335
rect 37274 57332 37280 57384
rect 37332 57372 37338 57384
rect 38105 57375 38163 57381
rect 38105 57372 38117 57375
rect 37332 57344 38117 57372
rect 37332 57332 37338 57344
rect 38105 57341 38117 57344
rect 38151 57372 38163 57375
rect 38286 57372 38292 57384
rect 38151 57344 38292 57372
rect 38151 57341 38163 57344
rect 38105 57335 38163 57341
rect 38286 57332 38292 57344
rect 38344 57332 38350 57384
rect 38381 57375 38439 57381
rect 38381 57341 38393 57375
rect 38427 57341 38439 57375
rect 38381 57335 38439 57341
rect 34480 57276 36492 57304
rect 34480 57264 34486 57276
rect 31202 57236 31208 57248
rect 28408 57208 29224 57236
rect 31163 57208 31208 57236
rect 28408 57196 28414 57208
rect 31202 57196 31208 57208
rect 31260 57196 31266 57248
rect 31573 57239 31631 57245
rect 31573 57205 31585 57239
rect 31619 57236 31631 57239
rect 32030 57236 32036 57248
rect 31619 57208 32036 57236
rect 31619 57205 31631 57208
rect 31573 57199 31631 57205
rect 32030 57196 32036 57208
rect 32088 57196 32094 57248
rect 33689 57239 33747 57245
rect 33689 57205 33701 57239
rect 33735 57236 33747 57239
rect 33870 57236 33876 57248
rect 33735 57208 33876 57236
rect 33735 57205 33747 57208
rect 33689 57199 33747 57205
rect 33870 57196 33876 57208
rect 33928 57196 33934 57248
rect 34606 57196 34612 57248
rect 34664 57236 34670 57248
rect 34793 57239 34851 57245
rect 34793 57236 34805 57239
rect 34664 57208 34805 57236
rect 34664 57196 34670 57208
rect 34793 57205 34805 57208
rect 34839 57205 34851 57239
rect 35342 57236 35348 57248
rect 35303 57208 35348 57236
rect 34793 57199 34851 57205
rect 35342 57196 35348 57208
rect 35400 57196 35406 57248
rect 37274 57196 37280 57248
rect 37332 57236 37338 57248
rect 38396 57236 38424 57335
rect 39942 57332 39948 57384
rect 40000 57372 40006 57384
rect 40313 57375 40371 57381
rect 40313 57372 40325 57375
rect 40000 57344 40325 57372
rect 40000 57332 40006 57344
rect 40313 57341 40325 57344
rect 40359 57341 40371 57375
rect 40313 57335 40371 57341
rect 40405 57375 40463 57381
rect 40405 57341 40417 57375
rect 40451 57341 40463 57375
rect 40405 57335 40463 57341
rect 40420 57304 40448 57335
rect 40494 57332 40500 57384
rect 40552 57372 40558 57384
rect 41432 57372 41460 57403
rect 42794 57400 42800 57452
rect 42852 57440 42858 57452
rect 43349 57443 43407 57449
rect 43349 57440 43361 57443
rect 42852 57412 43361 57440
rect 42852 57400 42858 57412
rect 43349 57409 43361 57412
rect 43395 57440 43407 57443
rect 43530 57440 43536 57452
rect 43395 57412 43536 57440
rect 43395 57409 43407 57412
rect 43349 57403 43407 57409
rect 43530 57400 43536 57412
rect 43588 57400 43594 57452
rect 44085 57443 44143 57449
rect 44085 57409 44097 57443
rect 44131 57440 44143 57443
rect 44910 57440 44916 57452
rect 44131 57412 44916 57440
rect 44131 57409 44143 57412
rect 44085 57403 44143 57409
rect 44910 57400 44916 57412
rect 44968 57400 44974 57452
rect 45554 57400 45560 57452
rect 45612 57440 45618 57452
rect 46017 57443 46075 57449
rect 46017 57440 46029 57443
rect 45612 57412 46029 57440
rect 45612 57400 45618 57412
rect 46017 57409 46029 57412
rect 46063 57440 46075 57443
rect 46382 57440 46388 57452
rect 46063 57412 46388 57440
rect 46063 57409 46075 57412
rect 46017 57403 46075 57409
rect 46382 57400 46388 57412
rect 46440 57400 46446 57452
rect 46750 57440 46756 57452
rect 46711 57412 46756 57440
rect 46750 57400 46756 57412
rect 46808 57400 46814 57452
rect 46934 57400 46940 57452
rect 46992 57440 46998 57452
rect 47578 57440 47584 57452
rect 46992 57412 47584 57440
rect 46992 57400 46998 57412
rect 47578 57400 47584 57412
rect 47636 57440 47642 57452
rect 47765 57443 47823 57449
rect 47765 57440 47777 57443
rect 47636 57412 47777 57440
rect 47636 57400 47642 57412
rect 47765 57409 47777 57412
rect 47811 57409 47823 57443
rect 47765 57403 47823 57409
rect 49694 57400 49700 57452
rect 49752 57440 49758 57452
rect 49789 57443 49847 57449
rect 49789 57440 49801 57443
rect 49752 57412 49801 57440
rect 49752 57400 49758 57412
rect 49789 57409 49801 57412
rect 49835 57409 49847 57443
rect 49789 57403 49847 57409
rect 51074 57400 51080 57452
rect 51132 57440 51138 57452
rect 51442 57440 51448 57452
rect 51132 57412 51448 57440
rect 51132 57400 51138 57412
rect 51442 57400 51448 57412
rect 51500 57440 51506 57452
rect 51629 57443 51687 57449
rect 51629 57440 51641 57443
rect 51500 57412 51641 57440
rect 51500 57400 51506 57412
rect 51629 57409 51641 57412
rect 51675 57409 51687 57443
rect 51629 57403 51687 57409
rect 53834 57400 53840 57452
rect 53892 57440 53898 57452
rect 53929 57443 53987 57449
rect 53929 57440 53941 57443
rect 53892 57412 53941 57440
rect 53892 57400 53898 57412
rect 53929 57409 53941 57412
rect 53975 57409 53987 57443
rect 53929 57403 53987 57409
rect 54294 57400 54300 57452
rect 54352 57440 54358 57452
rect 54665 57443 54723 57449
rect 54665 57440 54677 57443
rect 54352 57412 54677 57440
rect 54352 57400 54358 57412
rect 54665 57409 54677 57412
rect 54711 57409 54723 57443
rect 54665 57403 54723 57409
rect 55214 57400 55220 57452
rect 55272 57440 55278 57452
rect 55493 57443 55551 57449
rect 55493 57440 55505 57443
rect 55272 57412 55505 57440
rect 55272 57400 55278 57412
rect 55493 57409 55505 57412
rect 55539 57409 55551 57443
rect 55493 57403 55551 57409
rect 55674 57400 55680 57452
rect 55732 57440 55738 57452
rect 56229 57443 56287 57449
rect 56229 57440 56241 57443
rect 55732 57412 56241 57440
rect 55732 57400 55738 57412
rect 56229 57409 56241 57412
rect 56275 57409 56287 57443
rect 56229 57403 56287 57409
rect 43073 57375 43131 57381
rect 43073 57372 43085 57375
rect 40552 57344 40597 57372
rect 41432 57344 43085 57372
rect 40552 57332 40558 57344
rect 43073 57341 43085 57344
rect 43119 57372 43131 57375
rect 43990 57372 43996 57384
rect 43119 57344 43996 57372
rect 43119 57341 43131 57344
rect 43073 57335 43131 57341
rect 43990 57332 43996 57344
rect 44048 57332 44054 57384
rect 44361 57375 44419 57381
rect 44361 57341 44373 57375
rect 44407 57372 44419 57375
rect 44450 57372 44456 57384
rect 44407 57344 44456 57372
rect 44407 57341 44419 57344
rect 44361 57335 44419 57341
rect 44450 57332 44456 57344
rect 44508 57372 44514 57384
rect 50065 57375 50123 57381
rect 50065 57372 50077 57375
rect 44508 57344 50077 57372
rect 44508 57332 44514 57344
rect 50065 57341 50077 57344
rect 50111 57341 50123 57375
rect 50065 57335 50123 57341
rect 40954 57304 40960 57316
rect 40420 57276 40960 57304
rect 40954 57264 40960 57276
rect 41012 57264 41018 57316
rect 43162 57264 43168 57316
rect 43220 57304 43226 57316
rect 43220 57276 46060 57304
rect 43220 57264 43226 57276
rect 37332 57208 38424 57236
rect 37332 57196 37338 57208
rect 40126 57196 40132 57248
rect 40184 57236 40190 57248
rect 41049 57239 41107 57245
rect 41049 57236 41061 57239
rect 40184 57208 41061 57236
rect 40184 57196 40190 57208
rect 41049 57205 41061 57208
rect 41095 57205 41107 57239
rect 43898 57236 43904 57248
rect 43859 57208 43904 57236
rect 41049 57199 41107 57205
rect 43898 57196 43904 57208
rect 43956 57196 43962 57248
rect 44266 57236 44272 57248
rect 44227 57208 44272 57236
rect 44266 57196 44272 57208
rect 44324 57196 44330 57248
rect 44818 57236 44824 57248
rect 44779 57208 44824 57236
rect 44818 57196 44824 57208
rect 44876 57196 44882 57248
rect 45922 57236 45928 57248
rect 45883 57208 45928 57236
rect 45922 57196 45928 57208
rect 45980 57196 45986 57248
rect 46032 57236 46060 57276
rect 46382 57264 46388 57316
rect 46440 57304 46446 57316
rect 49053 57307 49111 57313
rect 49053 57304 49065 57307
rect 46440 57276 49065 57304
rect 46440 57264 46446 57276
rect 49053 57273 49065 57276
rect 49099 57273 49111 57307
rect 49053 57267 49111 57273
rect 49142 57264 49148 57316
rect 49200 57304 49206 57316
rect 51813 57307 51871 57313
rect 51813 57304 51825 57307
rect 49200 57276 51825 57304
rect 49200 57264 49206 57276
rect 51813 57273 51825 57276
rect 51859 57273 51871 57307
rect 51813 57267 51871 57273
rect 46569 57239 46627 57245
rect 46569 57236 46581 57239
rect 46032 57208 46581 57236
rect 46569 57205 46581 57208
rect 46615 57205 46627 57239
rect 54110 57236 54116 57248
rect 54071 57208 54116 57236
rect 46569 57199 46627 57205
rect 54110 57196 54116 57208
rect 54168 57196 54174 57248
rect 54202 57196 54208 57248
rect 54260 57236 54266 57248
rect 55677 57239 55735 57245
rect 55677 57236 55689 57239
rect 54260 57208 55689 57236
rect 54260 57196 54266 57208
rect 55677 57205 55689 57208
rect 55723 57205 55735 57239
rect 55677 57199 55735 57205
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 3694 57032 3700 57044
rect 3655 57004 3700 57032
rect 3694 56992 3700 57004
rect 3752 56992 3758 57044
rect 5994 56992 6000 57044
rect 6052 57032 6058 57044
rect 6089 57035 6147 57041
rect 6089 57032 6101 57035
rect 6052 57004 6101 57032
rect 6052 56992 6058 57004
rect 6089 57001 6101 57004
rect 6135 57001 6147 57035
rect 6089 56995 6147 57001
rect 7374 56992 7380 57044
rect 7432 57032 7438 57044
rect 7469 57035 7527 57041
rect 7469 57032 7481 57035
rect 7432 57004 7481 57032
rect 7432 56992 7438 57004
rect 7469 57001 7481 57004
rect 7515 57001 7527 57035
rect 7469 56995 7527 57001
rect 11514 56992 11520 57044
rect 11572 57032 11578 57044
rect 11609 57035 11667 57041
rect 11609 57032 11621 57035
rect 11572 57004 11621 57032
rect 11572 56992 11578 57004
rect 11609 57001 11621 57004
rect 11655 57001 11667 57035
rect 11609 56995 11667 57001
rect 12894 56992 12900 57044
rect 12952 57032 12958 57044
rect 12989 57035 13047 57041
rect 12989 57032 13001 57035
rect 12952 57004 13001 57032
rect 12952 56992 12958 57004
rect 12989 57001 13001 57004
rect 13035 57001 13047 57035
rect 12989 56995 13047 57001
rect 17034 56992 17040 57044
rect 17092 57032 17098 57044
rect 17129 57035 17187 57041
rect 17129 57032 17141 57035
rect 17092 57004 17141 57032
rect 17092 56992 17098 57004
rect 17129 57001 17141 57004
rect 17175 57001 17187 57035
rect 17129 56995 17187 57001
rect 18414 56992 18420 57044
rect 18472 57032 18478 57044
rect 19153 57035 19211 57041
rect 19153 57032 19165 57035
rect 18472 57004 19165 57032
rect 18472 56992 18478 57004
rect 19153 57001 19165 57004
rect 19199 57001 19211 57035
rect 19153 56995 19211 57001
rect 21174 56992 21180 57044
rect 21232 57032 21238 57044
rect 21269 57035 21327 57041
rect 21269 57032 21281 57035
rect 21232 57004 21281 57032
rect 21232 56992 21238 57004
rect 21269 57001 21281 57004
rect 21315 57001 21327 57035
rect 21269 56995 21327 57001
rect 23198 56992 23204 57044
rect 23256 57032 23262 57044
rect 24305 57035 24363 57041
rect 24305 57032 24317 57035
rect 23256 57004 24317 57032
rect 23256 56992 23262 57004
rect 24305 57001 24317 57004
rect 24351 57001 24363 57035
rect 25682 57032 25688 57044
rect 25643 57004 25688 57032
rect 24305 56995 24363 57001
rect 25682 56992 25688 57004
rect 25740 56992 25746 57044
rect 26970 56992 26976 57044
rect 27028 57032 27034 57044
rect 27157 57035 27215 57041
rect 27157 57032 27169 57035
rect 27028 57004 27169 57032
rect 27028 56992 27034 57004
rect 27157 57001 27169 57004
rect 27203 57001 27215 57035
rect 27157 56995 27215 57001
rect 28629 57035 28687 57041
rect 28629 57001 28641 57035
rect 28675 57032 28687 57035
rect 29822 57032 29828 57044
rect 28675 57004 29828 57032
rect 28675 57001 28687 57004
rect 28629 56995 28687 57001
rect 29822 56992 29828 57004
rect 29880 56992 29886 57044
rect 29917 57035 29975 57041
rect 29917 57001 29929 57035
rect 29963 57032 29975 57035
rect 30006 57032 30012 57044
rect 29963 57004 30012 57032
rect 29963 57001 29975 57004
rect 29917 56995 29975 57001
rect 30006 56992 30012 57004
rect 30064 56992 30070 57044
rect 30834 56992 30840 57044
rect 30892 57032 30898 57044
rect 31021 57035 31079 57041
rect 31021 57032 31033 57035
rect 30892 57004 31033 57032
rect 30892 56992 30898 57004
rect 31021 57001 31033 57004
rect 31067 57001 31079 57035
rect 31021 56995 31079 57001
rect 31386 56992 31392 57044
rect 31444 57032 31450 57044
rect 31665 57035 31723 57041
rect 31665 57032 31677 57035
rect 31444 57004 31677 57032
rect 31444 56992 31450 57004
rect 31665 57001 31677 57004
rect 31711 57001 31723 57035
rect 34238 57032 34244 57044
rect 34199 57004 34244 57032
rect 31665 56995 31723 57001
rect 34238 56992 34244 57004
rect 34296 56992 34302 57044
rect 34698 56992 34704 57044
rect 34756 57032 34762 57044
rect 35161 57035 35219 57041
rect 35161 57032 35173 57035
rect 34756 57004 35173 57032
rect 34756 56992 34762 57004
rect 35161 57001 35173 57004
rect 35207 57001 35219 57035
rect 35161 56995 35219 57001
rect 36722 56992 36728 57044
rect 36780 57032 36786 57044
rect 39850 57032 39856 57044
rect 36780 57004 39856 57032
rect 36780 56992 36786 57004
rect 39850 56992 39856 57004
rect 39908 56992 39914 57044
rect 41782 56992 41788 57044
rect 41840 57032 41846 57044
rect 43257 57035 43315 57041
rect 43257 57032 43269 57035
rect 41840 57004 43269 57032
rect 41840 56992 41846 57004
rect 43257 57001 43269 57004
rect 43303 57032 43315 57035
rect 44266 57032 44272 57044
rect 43303 57004 44272 57032
rect 43303 57001 43315 57004
rect 43257 56995 43315 57001
rect 44266 56992 44272 57004
rect 44324 56992 44330 57044
rect 46014 56992 46020 57044
rect 46072 57032 46078 57044
rect 47489 57035 47547 57041
rect 47489 57032 47501 57035
rect 46072 57004 47501 57032
rect 46072 56992 46078 57004
rect 47489 57001 47501 57004
rect 47535 57001 47547 57035
rect 47489 56995 47547 57001
rect 47854 56992 47860 57044
rect 47912 57032 47918 57044
rect 49697 57035 49755 57041
rect 49697 57032 49709 57035
rect 47912 57004 49709 57032
rect 47912 56992 47918 57004
rect 49697 57001 49709 57004
rect 49743 57001 49755 57035
rect 49697 56995 49755 57001
rect 50154 56992 50160 57044
rect 50212 57032 50218 57044
rect 50801 57035 50859 57041
rect 50801 57032 50813 57035
rect 50212 57004 50813 57032
rect 50212 56992 50218 57004
rect 50801 57001 50813 57004
rect 50847 57001 50859 57035
rect 50801 56995 50859 57001
rect 51534 56992 51540 57044
rect 51592 57032 51598 57044
rect 52089 57035 52147 57041
rect 52089 57032 52101 57035
rect 51592 57004 52101 57032
rect 51592 56992 51598 57004
rect 52089 57001 52101 57004
rect 52135 57001 52147 57035
rect 52089 56995 52147 57001
rect 52454 56992 52460 57044
rect 52512 57032 52518 57044
rect 52733 57035 52791 57041
rect 52733 57032 52745 57035
rect 52512 57004 52745 57032
rect 52512 56992 52518 57004
rect 52733 57001 52745 57004
rect 52779 57001 52791 57035
rect 52733 56995 52791 57001
rect 52914 56992 52920 57044
rect 52972 57032 52978 57044
rect 53377 57035 53435 57041
rect 53377 57032 53389 57035
rect 52972 57004 53389 57032
rect 52972 56992 52978 57004
rect 53377 57001 53389 57004
rect 53423 57001 53435 57035
rect 53377 56995 53435 57001
rect 53466 56992 53472 57044
rect 53524 57032 53530 57044
rect 54021 57035 54079 57041
rect 54021 57032 54033 57035
rect 53524 57004 54033 57032
rect 53524 56992 53530 57004
rect 54021 57001 54033 57004
rect 54067 57001 54079 57035
rect 54021 56995 54079 57001
rect 54754 56992 54760 57044
rect 54812 57032 54818 57044
rect 54849 57035 54907 57041
rect 54849 57032 54861 57035
rect 54812 57004 54861 57032
rect 54812 56992 54818 57004
rect 54849 57001 54861 57004
rect 54895 57001 54907 57035
rect 54849 56995 54907 57001
rect 55214 56992 55220 57044
rect 55272 57032 55278 57044
rect 55493 57035 55551 57041
rect 55493 57032 55505 57035
rect 55272 57004 55505 57032
rect 55272 56992 55278 57004
rect 55493 57001 55505 57004
rect 55539 57001 55551 57035
rect 55493 56995 55551 57001
rect 56134 56992 56140 57044
rect 56192 57032 56198 57044
rect 56229 57035 56287 57041
rect 56229 57032 56241 57035
rect 56192 57004 56241 57032
rect 56192 56992 56198 57004
rect 56229 57001 56241 57004
rect 56275 57001 56287 57035
rect 56229 56995 56287 57001
rect 19242 56924 19248 56976
rect 19300 56964 19306 56976
rect 22373 56967 22431 56973
rect 22373 56964 22385 56967
rect 19300 56936 22385 56964
rect 19300 56924 19306 56936
rect 22373 56933 22385 56936
rect 22419 56933 22431 56967
rect 22373 56927 22431 56933
rect 11330 56856 11336 56908
rect 11388 56896 11394 56908
rect 12345 56899 12403 56905
rect 12345 56896 12357 56899
rect 11388 56868 12357 56896
rect 11388 56856 11394 56868
rect 12345 56865 12357 56868
rect 12391 56896 12403 56899
rect 21358 56896 21364 56908
rect 12391 56868 21364 56896
rect 12391 56865 12403 56868
rect 12345 56859 12403 56865
rect 21358 56856 21364 56868
rect 21416 56856 21422 56908
rect 22388 56896 22416 56927
rect 22462 56924 22468 56976
rect 22520 56964 22526 56976
rect 27709 56967 27767 56973
rect 27709 56964 27721 56967
rect 22520 56936 27721 56964
rect 22520 56924 22526 56936
rect 27709 56933 27721 56936
rect 27755 56933 27767 56967
rect 27709 56927 27767 56933
rect 30282 56924 30288 56976
rect 30340 56964 30346 56976
rect 30469 56967 30527 56973
rect 30469 56964 30481 56967
rect 30340 56936 30481 56964
rect 30340 56924 30346 56936
rect 30469 56933 30481 56936
rect 30515 56964 30527 56967
rect 32217 56967 32275 56973
rect 32217 56964 32229 56967
rect 30515 56936 32229 56964
rect 30515 56933 30527 56936
rect 30469 56927 30527 56933
rect 32217 56933 32229 56936
rect 32263 56964 32275 56967
rect 32263 56936 33456 56964
rect 32263 56933 32275 56936
rect 32217 56927 32275 56933
rect 23661 56899 23719 56905
rect 23661 56896 23673 56899
rect 22388 56868 23673 56896
rect 23661 56865 23673 56868
rect 23707 56865 23719 56899
rect 23661 56859 23719 56865
rect 24026 56856 24032 56908
rect 24084 56896 24090 56908
rect 24854 56896 24860 56908
rect 24084 56868 24860 56896
rect 24084 56856 24090 56868
rect 24854 56856 24860 56868
rect 24912 56856 24918 56908
rect 25038 56896 25044 56908
rect 24999 56868 25044 56896
rect 25038 56856 25044 56868
rect 25096 56856 25102 56908
rect 25222 56856 25228 56908
rect 25280 56896 25286 56908
rect 27062 56896 27068 56908
rect 25280 56868 26924 56896
rect 27023 56868 27068 56896
rect 25280 56856 25286 56868
rect 22557 56831 22615 56837
rect 22557 56797 22569 56831
rect 22603 56828 22615 56831
rect 22646 56828 22652 56840
rect 22603 56800 22652 56828
rect 22603 56797 22615 56800
rect 22557 56791 22615 56797
rect 22646 56788 22652 56800
rect 22704 56788 22710 56840
rect 23750 56788 23756 56840
rect 23808 56828 23814 56840
rect 24210 56837 24216 56840
rect 24180 56831 24216 56837
rect 23808 56800 23853 56828
rect 23808 56788 23814 56800
rect 24180 56797 24192 56831
rect 24180 56791 24216 56797
rect 24210 56788 24216 56791
rect 24268 56788 24274 56840
rect 25130 56788 25136 56840
rect 25188 56828 25194 56840
rect 25590 56837 25596 56840
rect 25560 56831 25596 56837
rect 25188 56800 25233 56828
rect 25188 56788 25194 56800
rect 25560 56797 25572 56831
rect 25560 56791 25596 56797
rect 25590 56788 25596 56791
rect 25648 56788 25654 56840
rect 26326 56828 26332 56840
rect 26287 56800 26332 56828
rect 26326 56788 26332 56800
rect 26384 56788 26390 56840
rect 26418 56788 26424 56840
rect 26476 56828 26482 56840
rect 26896 56828 26924 56868
rect 27062 56856 27068 56868
rect 27120 56856 27126 56908
rect 27614 56896 27620 56908
rect 27172 56868 27620 56896
rect 27172 56828 27200 56868
rect 27614 56856 27620 56868
rect 27672 56896 27678 56908
rect 27672 56868 27752 56896
rect 27672 56856 27678 56868
rect 26476 56800 26521 56828
rect 26896 56800 27200 56828
rect 26476 56788 26482 56800
rect 27522 56788 27528 56840
rect 27580 56828 27586 56840
rect 27724 56828 27752 56868
rect 27798 56856 27804 56908
rect 27856 56896 27862 56908
rect 27856 56868 28488 56896
rect 27856 56856 27862 56868
rect 27982 56828 27988 56840
rect 27580 56800 27625 56828
rect 27724 56800 27988 56828
rect 27580 56788 27586 56800
rect 27982 56788 27988 56800
rect 28040 56828 28046 56840
rect 28460 56837 28488 56868
rect 28534 56856 28540 56908
rect 28592 56896 28598 56908
rect 29457 56899 29515 56905
rect 29457 56896 29469 56899
rect 28592 56868 29469 56896
rect 28592 56856 28598 56868
rect 29457 56865 29469 56868
rect 29503 56896 29515 56899
rect 33042 56896 33048 56908
rect 29503 56868 33048 56896
rect 29503 56865 29515 56868
rect 29457 56859 29515 56865
rect 33042 56856 33048 56868
rect 33100 56856 33106 56908
rect 33428 56896 33456 56936
rect 33686 56924 33692 56976
rect 33744 56964 33750 56976
rect 36081 56967 36139 56973
rect 36081 56964 36093 56967
rect 33744 56936 36093 56964
rect 33744 56924 33750 56936
rect 36081 56933 36093 56936
rect 36127 56933 36139 56967
rect 36081 56927 36139 56933
rect 36262 56924 36268 56976
rect 36320 56964 36326 56976
rect 41138 56964 41144 56976
rect 36320 56936 41144 56964
rect 36320 56924 36326 56936
rect 41138 56924 41144 56936
rect 41196 56924 41202 56976
rect 43346 56964 43352 56976
rect 41800 56936 43352 56964
rect 33870 56896 33876 56908
rect 33428 56868 33876 56896
rect 28353 56831 28411 56837
rect 28353 56828 28365 56831
rect 28040 56800 28365 56828
rect 28040 56788 28046 56800
rect 28353 56797 28365 56800
rect 28399 56797 28411 56831
rect 28353 56791 28411 56797
rect 28445 56831 28503 56837
rect 28445 56797 28457 56831
rect 28491 56797 28503 56831
rect 28718 56828 28724 56840
rect 28679 56800 28724 56828
rect 28445 56791 28503 56797
rect 28718 56788 28724 56800
rect 28776 56788 28782 56840
rect 28810 56788 28816 56840
rect 28868 56828 28874 56840
rect 29181 56831 29239 56837
rect 29181 56828 29193 56831
rect 28868 56800 29193 56828
rect 28868 56788 28874 56800
rect 29181 56797 29193 56800
rect 29227 56797 29239 56831
rect 29365 56831 29423 56837
rect 29365 56828 29377 56831
rect 29181 56791 29239 56797
rect 29288 56800 29377 56828
rect 7282 56720 7288 56772
rect 7340 56760 7346 56772
rect 28169 56763 28227 56769
rect 28169 56760 28181 56763
rect 7340 56732 26280 56760
rect 7340 56720 7346 56732
rect 16942 56652 16948 56704
rect 17000 56692 17006 56704
rect 23109 56695 23167 56701
rect 23109 56692 23121 56695
rect 17000 56664 23121 56692
rect 17000 56652 17006 56664
rect 23109 56661 23121 56664
rect 23155 56692 23167 56695
rect 24026 56692 24032 56704
rect 23155 56664 24032 56692
rect 23155 56661 23167 56664
rect 23109 56655 23167 56661
rect 24026 56652 24032 56664
rect 24084 56652 24090 56704
rect 24121 56695 24179 56701
rect 24121 56661 24133 56695
rect 24167 56692 24179 56695
rect 24762 56692 24768 56704
rect 24167 56664 24768 56692
rect 24167 56661 24179 56664
rect 24121 56655 24179 56661
rect 24762 56652 24768 56664
rect 24820 56652 24826 56704
rect 25501 56695 25559 56701
rect 25501 56661 25513 56695
rect 25547 56692 25559 56695
rect 25682 56692 25688 56704
rect 25547 56664 25688 56692
rect 25547 56661 25559 56664
rect 25501 56655 25559 56661
rect 25682 56652 25688 56664
rect 25740 56652 25746 56704
rect 26142 56692 26148 56704
rect 26103 56664 26148 56692
rect 26142 56652 26148 56664
rect 26200 56652 26206 56704
rect 26252 56692 26280 56732
rect 26436 56732 28181 56760
rect 26436 56692 26464 56732
rect 28169 56729 28181 56732
rect 28215 56729 28227 56763
rect 28169 56723 28227 56729
rect 28626 56720 28632 56772
rect 28684 56760 28690 56772
rect 28902 56760 28908 56772
rect 28684 56732 28908 56760
rect 28684 56720 28690 56732
rect 28902 56720 28908 56732
rect 28960 56760 28966 56772
rect 29288 56760 29316 56800
rect 29365 56797 29377 56800
rect 29411 56797 29423 56831
rect 29365 56791 29423 56797
rect 29546 56788 29552 56840
rect 29604 56828 29610 56840
rect 29730 56828 29736 56840
rect 29604 56800 29649 56828
rect 29691 56800 29736 56828
rect 29604 56788 29610 56800
rect 29730 56788 29736 56800
rect 29788 56788 29794 56840
rect 31662 56788 31668 56840
rect 31720 56828 31726 56840
rect 31790 56831 31848 56837
rect 31790 56828 31802 56831
rect 31720 56800 31802 56828
rect 31720 56788 31726 56800
rect 31790 56797 31802 56800
rect 31836 56797 31848 56831
rect 32306 56828 32312 56840
rect 32267 56800 32312 56828
rect 31790 56791 31848 56797
rect 32306 56788 32312 56800
rect 32364 56788 32370 56840
rect 33428 56837 33456 56868
rect 33870 56856 33876 56868
rect 33928 56856 33934 56908
rect 35618 56896 35624 56908
rect 35531 56868 35624 56896
rect 33413 56831 33471 56837
rect 33413 56797 33425 56831
rect 33459 56797 33471 56831
rect 33413 56791 33471 56797
rect 33505 56831 33563 56837
rect 33505 56797 33517 56831
rect 33551 56797 33563 56831
rect 33686 56828 33692 56840
rect 33647 56800 33692 56828
rect 33505 56791 33563 56797
rect 28960 56732 29316 56760
rect 33512 56760 33540 56791
rect 33686 56788 33692 56800
rect 33744 56788 33750 56840
rect 33778 56788 33784 56840
rect 33836 56828 33842 56840
rect 35544 56837 35572 56868
rect 35618 56856 35624 56868
rect 35676 56896 35682 56908
rect 37829 56899 37887 56905
rect 37829 56896 37841 56899
rect 35676 56868 37841 56896
rect 35676 56856 35682 56868
rect 37829 56865 37841 56868
rect 37875 56865 37887 56899
rect 37829 56859 37887 56865
rect 38197 56899 38255 56905
rect 38197 56865 38209 56899
rect 38243 56896 38255 56899
rect 38378 56896 38384 56908
rect 38243 56868 38384 56896
rect 38243 56865 38255 56868
rect 38197 56859 38255 56865
rect 38378 56856 38384 56868
rect 38436 56856 38442 56908
rect 38654 56856 38660 56908
rect 38712 56896 38718 56908
rect 38933 56899 38991 56905
rect 38933 56896 38945 56899
rect 38712 56868 38945 56896
rect 38712 56856 38718 56868
rect 38933 56865 38945 56868
rect 38979 56865 38991 56899
rect 38933 56859 38991 56865
rect 40589 56899 40647 56905
rect 40589 56865 40601 56899
rect 40635 56896 40647 56899
rect 41230 56896 41236 56908
rect 40635 56868 41236 56896
rect 40635 56865 40647 56868
rect 40589 56859 40647 56865
rect 41230 56856 41236 56868
rect 41288 56896 41294 56908
rect 41800 56896 41828 56936
rect 43346 56924 43352 56936
rect 43404 56924 43410 56976
rect 43714 56924 43720 56976
rect 43772 56964 43778 56976
rect 46845 56967 46903 56973
rect 46845 56964 46857 56967
rect 43772 56936 46857 56964
rect 43772 56924 43778 56936
rect 46845 56933 46857 56936
rect 46891 56933 46903 56967
rect 46845 56927 46903 56933
rect 50614 56924 50620 56976
rect 50672 56964 50678 56976
rect 51445 56967 51503 56973
rect 51445 56964 51457 56967
rect 50672 56936 51457 56964
rect 50672 56924 50678 56936
rect 51445 56933 51457 56936
rect 51491 56933 51503 56967
rect 51445 56927 51503 56933
rect 43898 56896 43904 56908
rect 41288 56868 41644 56896
rect 41800 56868 41920 56896
rect 43859 56868 43904 56896
rect 41288 56856 41294 56868
rect 35529 56831 35587 56837
rect 33836 56800 33881 56828
rect 33836 56788 33842 56800
rect 35529 56797 35541 56831
rect 35575 56797 35587 56831
rect 35986 56828 35992 56840
rect 35947 56800 35992 56828
rect 35529 56791 35587 56797
rect 35986 56788 35992 56800
rect 36044 56788 36050 56840
rect 36262 56828 36268 56840
rect 36223 56800 36268 56828
rect 36262 56788 36268 56800
rect 36320 56788 36326 56840
rect 36541 56831 36599 56837
rect 36541 56797 36553 56831
rect 36587 56828 36599 56831
rect 36630 56828 36636 56840
rect 36587 56800 36636 56828
rect 36587 56797 36599 56800
rect 36541 56791 36599 56797
rect 36630 56788 36636 56800
rect 36688 56788 36694 56840
rect 36814 56828 36820 56840
rect 36775 56800 36820 56828
rect 36814 56788 36820 56800
rect 36872 56788 36878 56840
rect 37369 56831 37427 56837
rect 37369 56797 37381 56831
rect 37415 56828 37427 56831
rect 37550 56828 37556 56840
rect 37415 56800 37556 56828
rect 37415 56797 37427 56800
rect 37369 56791 37427 56797
rect 37550 56788 37556 56800
rect 37608 56788 37614 56840
rect 38010 56828 38016 56840
rect 37971 56800 38016 56828
rect 38010 56788 38016 56800
rect 38068 56788 38074 56840
rect 38102 56788 38108 56840
rect 38160 56828 38166 56840
rect 38289 56831 38347 56837
rect 38160 56800 38205 56828
rect 38160 56788 38166 56800
rect 38289 56797 38301 56831
rect 38335 56828 38347 56831
rect 38746 56828 38752 56840
rect 38335 56800 38752 56828
rect 38335 56797 38347 56800
rect 38289 56791 38347 56797
rect 38746 56788 38752 56800
rect 38804 56788 38810 56840
rect 39022 56788 39028 56840
rect 39080 56828 39086 56840
rect 39209 56831 39267 56837
rect 39209 56828 39221 56831
rect 39080 56800 39221 56828
rect 39080 56788 39086 56800
rect 39209 56797 39221 56800
rect 39255 56797 39267 56831
rect 39209 56791 39267 56797
rect 39850 56788 39856 56840
rect 39908 56828 39914 56840
rect 40497 56831 40555 56837
rect 40497 56828 40509 56831
rect 39908 56800 40509 56828
rect 39908 56788 39914 56800
rect 40497 56797 40509 56800
rect 40543 56828 40555 56831
rect 40770 56828 40776 56840
rect 40543 56800 40776 56828
rect 40543 56797 40555 56800
rect 40497 56791 40555 56797
rect 40770 56788 40776 56800
rect 40828 56788 40834 56840
rect 40954 56828 40960 56840
rect 40926 56800 40960 56828
rect 40954 56788 40960 56800
rect 41012 56837 41018 56840
rect 41012 56831 41074 56837
rect 41012 56797 41028 56831
rect 41062 56828 41074 56831
rect 41506 56828 41512 56840
rect 41062 56800 41512 56828
rect 41062 56797 41074 56800
rect 41012 56791 41074 56797
rect 41012 56788 41018 56791
rect 41506 56788 41512 56800
rect 41564 56788 41570 56840
rect 41616 56828 41644 56868
rect 41782 56828 41788 56840
rect 41616 56800 41788 56828
rect 41782 56788 41788 56800
rect 41840 56788 41846 56840
rect 41892 56837 41920 56868
rect 43898 56856 43904 56868
rect 43956 56856 43962 56908
rect 48314 56856 48320 56908
rect 48372 56896 48378 56908
rect 48409 56899 48467 56905
rect 48409 56896 48421 56899
rect 48372 56868 48421 56896
rect 48372 56856 48378 56868
rect 48409 56865 48421 56868
rect 48455 56865 48467 56899
rect 48409 56859 48467 56865
rect 41877 56831 41935 56837
rect 41877 56797 41889 56831
rect 41923 56797 41935 56831
rect 41877 56791 41935 56797
rect 41966 56788 41972 56840
rect 42024 56806 42030 56840
rect 42073 56831 42131 56837
rect 42073 56806 42085 56831
rect 42024 56797 42085 56806
rect 42119 56797 42131 56831
rect 42024 56791 42131 56797
rect 42163 56831 42221 56837
rect 42163 56797 42175 56831
rect 42209 56828 42221 56831
rect 42889 56831 42947 56837
rect 42889 56828 42901 56831
rect 42209 56800 42901 56828
rect 42209 56797 42221 56800
rect 42163 56791 42221 56797
rect 42889 56797 42901 56800
rect 42935 56797 42947 56831
rect 42889 56791 42947 56797
rect 43073 56831 43131 56837
rect 43073 56797 43085 56831
rect 43119 56828 43131 56831
rect 43162 56828 43168 56840
rect 43119 56800 43168 56828
rect 43119 56797 43131 56800
rect 43073 56791 43131 56797
rect 42024 56788 42124 56791
rect 43162 56788 43168 56800
rect 43220 56788 43226 56840
rect 43346 56828 43352 56840
rect 43307 56800 43352 56828
rect 43346 56788 43352 56800
rect 43404 56828 43410 56840
rect 43622 56828 43628 56840
rect 43404 56800 43628 56828
rect 43404 56788 43410 56800
rect 43622 56788 43628 56800
rect 43680 56788 43686 56840
rect 44082 56828 44088 56840
rect 44043 56800 44088 56828
rect 44082 56788 44088 56800
rect 44140 56788 44146 56840
rect 44450 56828 44456 56840
rect 44411 56800 44456 56828
rect 44450 56788 44456 56800
rect 44508 56788 44514 56840
rect 44729 56831 44787 56837
rect 44729 56797 44741 56831
rect 44775 56797 44787 56831
rect 45186 56828 45192 56840
rect 45147 56800 45192 56828
rect 44729 56791 44787 56797
rect 41984 56778 42124 56788
rect 34422 56760 34428 56772
rect 33512 56732 34428 56760
rect 28960 56720 28966 56732
rect 34422 56720 34428 56732
rect 34480 56720 34486 56772
rect 35345 56763 35403 56769
rect 35345 56729 35357 56763
rect 35391 56760 35403 56763
rect 35802 56760 35808 56772
rect 35391 56732 35808 56760
rect 35391 56729 35403 56732
rect 35345 56723 35403 56729
rect 35802 56720 35808 56732
rect 35860 56720 35866 56772
rect 42242 56720 42248 56772
rect 42300 56760 42306 56772
rect 43993 56763 44051 56769
rect 43993 56760 44005 56763
rect 42300 56732 44005 56760
rect 42300 56720 42306 56732
rect 43993 56729 44005 56732
rect 44039 56729 44051 56763
rect 44744 56760 44772 56791
rect 45186 56788 45192 56800
rect 45244 56788 45250 56840
rect 45830 56828 45836 56840
rect 45791 56800 45836 56828
rect 45830 56788 45836 56800
rect 45888 56788 45894 56840
rect 48682 56828 48688 56840
rect 48643 56800 48688 56828
rect 48682 56788 48688 56800
rect 48740 56788 48746 56840
rect 45002 56760 45008 56772
rect 44744 56732 45008 56760
rect 43993 56723 44051 56729
rect 45002 56720 45008 56732
rect 45060 56760 45066 56772
rect 54110 56760 54116 56772
rect 45060 56732 54116 56760
rect 45060 56720 45066 56732
rect 54110 56720 54116 56732
rect 54168 56720 54174 56772
rect 26252 56664 26464 56692
rect 26510 56652 26516 56704
rect 26568 56692 26574 56704
rect 27525 56695 27583 56701
rect 27525 56692 27537 56695
rect 26568 56664 27537 56692
rect 26568 56652 26574 56664
rect 27525 56661 27537 56664
rect 27571 56692 27583 56695
rect 29546 56692 29552 56704
rect 27571 56664 29552 56692
rect 27571 56661 27583 56664
rect 27525 56655 27583 56661
rect 29546 56652 29552 56664
rect 29604 56652 29610 56704
rect 30834 56652 30840 56704
rect 30892 56692 30898 56704
rect 31849 56695 31907 56701
rect 31849 56692 31861 56695
rect 30892 56664 31861 56692
rect 30892 56652 30898 56664
rect 31849 56661 31861 56664
rect 31895 56692 31907 56695
rect 32030 56692 32036 56704
rect 31895 56664 32036 56692
rect 31895 56661 31907 56664
rect 31849 56655 31907 56661
rect 32030 56652 32036 56664
rect 32088 56652 32094 56704
rect 33226 56692 33232 56704
rect 33187 56664 33232 56692
rect 33226 56652 33232 56664
rect 33284 56652 33290 56704
rect 34514 56652 34520 56704
rect 34572 56692 34578 56704
rect 39482 56692 39488 56704
rect 34572 56664 39488 56692
rect 34572 56652 34578 56664
rect 39482 56652 39488 56664
rect 39540 56652 39546 56704
rect 40954 56692 40960 56704
rect 40915 56664 40960 56692
rect 40954 56652 40960 56664
rect 41012 56652 41018 56704
rect 41138 56692 41144 56704
rect 41099 56664 41144 56692
rect 41138 56652 41144 56664
rect 41196 56652 41202 56704
rect 41601 56695 41659 56701
rect 41601 56661 41613 56695
rect 41647 56692 41659 56695
rect 41966 56692 41972 56704
rect 41647 56664 41972 56692
rect 41647 56661 41659 56664
rect 41601 56655 41659 56661
rect 41966 56652 41972 56664
rect 42024 56652 42030 56704
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 23569 56491 23627 56497
rect 23569 56457 23581 56491
rect 23615 56488 23627 56491
rect 23750 56488 23756 56500
rect 23615 56460 23756 56488
rect 23615 56457 23627 56460
rect 23569 56451 23627 56457
rect 23750 56448 23756 56460
rect 23808 56448 23814 56500
rect 25590 56488 25596 56500
rect 25424 56460 25596 56488
rect 22554 56312 22560 56364
rect 22612 56352 22618 56364
rect 22649 56355 22707 56361
rect 22649 56352 22661 56355
rect 22612 56324 22661 56352
rect 22612 56312 22618 56324
rect 22649 56321 22661 56324
rect 22695 56321 22707 56355
rect 22649 56315 22707 56321
rect 23385 56355 23443 56361
rect 23385 56321 23397 56355
rect 23431 56352 23443 56355
rect 24029 56355 24087 56361
rect 24029 56352 24041 56355
rect 23431 56324 24041 56352
rect 23431 56321 23443 56324
rect 23385 56315 23443 56321
rect 24029 56321 24041 56324
rect 24075 56321 24087 56355
rect 24029 56315 24087 56321
rect 24210 56312 24216 56364
rect 24268 56352 24274 56364
rect 25424 56361 25452 56460
rect 25590 56448 25596 56460
rect 25648 56488 25654 56500
rect 28445 56491 28503 56497
rect 25648 56460 28396 56488
rect 25648 56448 25654 56460
rect 26234 56380 26240 56432
rect 26292 56420 26298 56432
rect 26329 56423 26387 56429
rect 26329 56420 26341 56423
rect 26292 56392 26341 56420
rect 26292 56380 26298 56392
rect 26329 56389 26341 56392
rect 26375 56420 26387 56423
rect 26375 56392 27384 56420
rect 26375 56389 26387 56392
rect 26329 56383 26387 56389
rect 25409 56355 25467 56361
rect 24268 56324 24361 56352
rect 24268 56312 24274 56324
rect 25409 56321 25421 56355
rect 25455 56321 25467 56355
rect 25866 56352 25872 56364
rect 25409 56315 25467 56321
rect 25516 56324 25872 56352
rect 24228 56216 24256 56312
rect 24397 56287 24455 56293
rect 24397 56253 24409 56287
rect 24443 56284 24455 56287
rect 24486 56284 24492 56296
rect 24443 56256 24492 56284
rect 24443 56253 24455 56256
rect 24397 56247 24455 56253
rect 24486 56244 24492 56256
rect 24544 56244 24550 56296
rect 24854 56244 24860 56296
rect 24912 56284 24918 56296
rect 25516 56284 25544 56324
rect 25866 56312 25872 56324
rect 25924 56352 25930 56364
rect 26053 56355 26111 56361
rect 26053 56352 26065 56355
rect 25924 56324 26065 56352
rect 25924 56312 25930 56324
rect 26053 56321 26065 56324
rect 26099 56352 26111 56355
rect 26418 56352 26424 56364
rect 26099 56324 26424 56352
rect 26099 56321 26111 56324
rect 26053 56315 26111 56321
rect 26418 56312 26424 56324
rect 26476 56312 26482 56364
rect 24912 56256 25544 56284
rect 25593 56287 25651 56293
rect 24912 56244 24918 56256
rect 25593 56253 25605 56287
rect 25639 56284 25651 56287
rect 26528 56284 26556 56392
rect 27157 56355 27215 56361
rect 27157 56321 27169 56355
rect 27203 56321 27215 56355
rect 27157 56315 27215 56321
rect 27356 56352 27384 56392
rect 27890 56380 27896 56432
rect 27948 56420 27954 56432
rect 28077 56423 28135 56429
rect 28077 56420 28089 56423
rect 27948 56392 28089 56420
rect 27948 56380 27954 56392
rect 28077 56389 28089 56392
rect 28123 56389 28135 56423
rect 28258 56420 28264 56432
rect 28219 56392 28264 56420
rect 28077 56383 28135 56389
rect 28258 56380 28264 56392
rect 28316 56380 28322 56432
rect 28368 56420 28396 56460
rect 28445 56457 28457 56491
rect 28491 56488 28503 56491
rect 28718 56488 28724 56500
rect 28491 56460 28724 56488
rect 28491 56457 28503 56460
rect 28445 56451 28503 56457
rect 28718 56448 28724 56460
rect 28776 56448 28782 56500
rect 28902 56448 28908 56500
rect 28960 56488 28966 56500
rect 32033 56491 32091 56497
rect 32033 56488 32045 56491
rect 28960 56460 32045 56488
rect 28960 56448 28966 56460
rect 32033 56457 32045 56460
rect 32079 56457 32091 56491
rect 32033 56451 32091 56457
rect 32214 56448 32220 56500
rect 32272 56488 32278 56500
rect 32272 56460 33732 56488
rect 32272 56448 32278 56460
rect 33045 56423 33103 56429
rect 33045 56420 33057 56423
rect 28368 56392 33057 56420
rect 33045 56389 33057 56392
rect 33091 56389 33103 56423
rect 33704 56420 33732 56460
rect 33778 56448 33784 56500
rect 33836 56488 33842 56500
rect 33965 56491 34023 56497
rect 33965 56488 33977 56491
rect 33836 56460 33977 56488
rect 33836 56448 33842 56460
rect 33965 56457 33977 56460
rect 34011 56457 34023 56491
rect 35526 56488 35532 56500
rect 35487 56460 35532 56488
rect 33965 56451 34023 56457
rect 35526 56448 35532 56460
rect 35584 56448 35590 56500
rect 36814 56448 36820 56500
rect 36872 56488 36878 56500
rect 37001 56491 37059 56497
rect 37001 56488 37013 56491
rect 36872 56460 37013 56488
rect 36872 56448 36878 56460
rect 37001 56457 37013 56460
rect 37047 56457 37059 56491
rect 37001 56451 37059 56457
rect 39482 56448 39488 56500
rect 39540 56488 39546 56500
rect 39577 56491 39635 56497
rect 39577 56488 39589 56491
rect 39540 56460 39589 56488
rect 39540 56448 39546 56460
rect 39577 56457 39589 56460
rect 39623 56457 39635 56491
rect 40126 56488 40132 56500
rect 39577 56451 39635 56457
rect 39776 56460 40132 56488
rect 35342 56420 35348 56432
rect 33704 56392 35348 56420
rect 33045 56383 33103 56389
rect 35342 56380 35348 56392
rect 35400 56380 35406 56432
rect 37458 56420 37464 56432
rect 35452 56392 37464 56420
rect 28810 56352 28816 56364
rect 27356 56324 28816 56352
rect 25639 56256 26556 56284
rect 25639 56253 25651 56256
rect 25593 56247 25651 56253
rect 27172 56216 27200 56315
rect 27356 56296 27384 56324
rect 28810 56312 28816 56324
rect 28868 56312 28874 56364
rect 28994 56312 29000 56364
rect 29052 56352 29058 56364
rect 29641 56355 29699 56361
rect 29641 56352 29653 56355
rect 29052 56324 29653 56352
rect 29052 56312 29058 56324
rect 29641 56321 29653 56324
rect 29687 56321 29699 56355
rect 29641 56315 29699 56321
rect 31113 56355 31171 56361
rect 31113 56321 31125 56355
rect 31159 56350 31171 56355
rect 31662 56352 31668 56364
rect 31312 56350 31668 56352
rect 31159 56324 31668 56350
rect 31159 56322 31340 56324
rect 31159 56321 31171 56322
rect 31113 56315 31171 56321
rect 31662 56312 31668 56324
rect 31720 56312 31726 56364
rect 32214 56312 32220 56364
rect 32272 56352 32278 56364
rect 33226 56352 33232 56364
rect 32272 56324 32904 56352
rect 33187 56324 33232 56352
rect 32272 56312 32278 56324
rect 27338 56284 27344 56296
rect 27299 56256 27344 56284
rect 27338 56244 27344 56256
rect 27396 56244 27402 56296
rect 27982 56244 27988 56296
rect 28040 56284 28046 56296
rect 29822 56284 29828 56296
rect 28040 56256 29828 56284
rect 28040 56244 28046 56256
rect 29822 56244 29828 56256
rect 29880 56244 29886 56296
rect 30834 56244 30840 56296
rect 30892 56284 30898 56296
rect 30929 56287 30987 56293
rect 30929 56284 30941 56287
rect 30892 56256 30941 56284
rect 30892 56244 30898 56256
rect 30929 56253 30941 56256
rect 30975 56253 30987 56287
rect 30929 56247 30987 56253
rect 31021 56287 31079 56293
rect 31021 56253 31033 56287
rect 31067 56253 31079 56287
rect 31021 56247 31079 56253
rect 31205 56287 31263 56293
rect 31205 56253 31217 56287
rect 31251 56253 31263 56287
rect 31205 56247 31263 56253
rect 32493 56287 32551 56293
rect 32493 56253 32505 56287
rect 32539 56284 32551 56287
rect 32766 56284 32772 56296
rect 32539 56256 32772 56284
rect 32539 56253 32551 56256
rect 32493 56247 32551 56253
rect 27522 56216 27528 56228
rect 24228 56188 27108 56216
rect 27172 56188 27528 56216
rect 24578 56108 24584 56160
rect 24636 56148 24642 56160
rect 25225 56151 25283 56157
rect 25225 56148 25237 56151
rect 24636 56120 25237 56148
rect 24636 56108 24642 56120
rect 25225 56117 25237 56120
rect 25271 56117 25283 56151
rect 25225 56111 25283 56117
rect 26602 56108 26608 56160
rect 26660 56148 26666 56160
rect 26973 56151 27031 56157
rect 26973 56148 26985 56151
rect 26660 56120 26985 56148
rect 26660 56108 26666 56120
rect 26973 56117 26985 56120
rect 27019 56117 27031 56151
rect 27080 56148 27108 56188
rect 27522 56176 27528 56188
rect 27580 56216 27586 56228
rect 28718 56216 28724 56228
rect 27580 56188 28724 56216
rect 27580 56176 27586 56188
rect 28718 56176 28724 56188
rect 28776 56176 28782 56228
rect 28828 56188 29592 56216
rect 28828 56148 28856 56188
rect 27080 56120 28856 56148
rect 26973 56111 27031 56117
rect 29362 56108 29368 56160
rect 29420 56148 29426 56160
rect 29457 56151 29515 56157
rect 29457 56148 29469 56151
rect 29420 56120 29469 56148
rect 29420 56108 29426 56120
rect 29457 56117 29469 56120
rect 29503 56117 29515 56151
rect 29564 56148 29592 56188
rect 29730 56176 29736 56228
rect 29788 56216 29794 56228
rect 31036 56216 31064 56247
rect 31110 56216 31116 56228
rect 29788 56188 31116 56216
rect 29788 56176 29794 56188
rect 31110 56176 31116 56188
rect 31168 56176 31174 56228
rect 31220 56160 31248 56247
rect 32766 56244 32772 56256
rect 32824 56244 32830 56296
rect 32876 56284 32904 56324
rect 33226 56312 33232 56324
rect 33284 56312 33290 56364
rect 34146 56352 34152 56364
rect 34107 56324 34152 56352
rect 34146 56312 34152 56324
rect 34204 56312 34210 56364
rect 34422 56312 34428 56364
rect 34480 56352 34486 56364
rect 35452 56352 35480 56392
rect 37458 56380 37464 56392
rect 37516 56380 37522 56432
rect 38194 56380 38200 56432
rect 38252 56420 38258 56432
rect 38838 56420 38844 56432
rect 38252 56392 38844 56420
rect 38252 56380 38258 56392
rect 38838 56380 38844 56392
rect 38896 56380 38902 56432
rect 35618 56352 35624 56364
rect 34480 56324 34525 56352
rect 34624 56324 35480 56352
rect 35579 56324 35624 56352
rect 34480 56312 34486 56324
rect 33318 56284 33324 56296
rect 32876 56256 33324 56284
rect 33318 56244 33324 56256
rect 33376 56244 33382 56296
rect 33505 56287 33563 56293
rect 33505 56253 33517 56287
rect 33551 56253 33563 56287
rect 33505 56247 33563 56253
rect 30745 56151 30803 56157
rect 30745 56148 30757 56151
rect 29564 56120 30757 56148
rect 29457 56111 29515 56117
rect 30745 56117 30757 56120
rect 30791 56117 30803 56151
rect 30745 56111 30803 56117
rect 31202 56108 31208 56160
rect 31260 56108 31266 56160
rect 32401 56151 32459 56157
rect 32401 56117 32413 56151
rect 32447 56148 32459 56151
rect 32490 56148 32496 56160
rect 32447 56120 32496 56148
rect 32447 56117 32459 56120
rect 32401 56111 32459 56117
rect 32490 56108 32496 56120
rect 32548 56108 32554 56160
rect 33410 56148 33416 56160
rect 33371 56120 33416 56148
rect 33410 56108 33416 56120
rect 33468 56108 33474 56160
rect 33520 56148 33548 56247
rect 33870 56244 33876 56296
rect 33928 56284 33934 56296
rect 34330 56284 34336 56296
rect 33928 56256 34336 56284
rect 33928 56244 33934 56256
rect 34330 56244 34336 56256
rect 34388 56284 34394 56296
rect 34624 56284 34652 56324
rect 35618 56312 35624 56324
rect 35676 56312 35682 56364
rect 35802 56352 35808 56364
rect 35763 56324 35808 56352
rect 35802 56312 35808 56324
rect 35860 56312 35866 56364
rect 35986 56352 35992 56364
rect 35947 56324 35992 56352
rect 35986 56312 35992 56324
rect 36044 56352 36050 56364
rect 36446 56352 36452 56364
rect 36044 56324 36452 56352
rect 36044 56312 36050 56324
rect 36446 56312 36452 56324
rect 36504 56312 36510 56364
rect 37369 56355 37427 56361
rect 37369 56321 37381 56355
rect 37415 56352 37427 56355
rect 37918 56352 37924 56364
rect 37415 56324 37924 56352
rect 37415 56321 37427 56324
rect 37369 56315 37427 56321
rect 37918 56312 37924 56324
rect 37976 56312 37982 56364
rect 39776 56361 39804 56460
rect 40126 56448 40132 56460
rect 40184 56448 40190 56500
rect 40494 56448 40500 56500
rect 40552 56488 40558 56500
rect 40957 56491 41015 56497
rect 40957 56488 40969 56491
rect 40552 56460 40969 56488
rect 40552 56448 40558 56460
rect 40957 56457 40969 56460
rect 41003 56457 41015 56491
rect 40957 56451 41015 56457
rect 41874 56448 41880 56500
rect 41932 56488 41938 56500
rect 42886 56488 42892 56500
rect 41932 56460 42892 56488
rect 41932 56448 41938 56460
rect 42886 56448 42892 56460
rect 42944 56448 42950 56500
rect 44266 56488 44272 56500
rect 44179 56460 44272 56488
rect 44266 56448 44272 56460
rect 44324 56488 44330 56500
rect 45002 56488 45008 56500
rect 44324 56460 45008 56488
rect 44324 56448 44330 56460
rect 45002 56448 45008 56460
rect 45060 56448 45066 56500
rect 49694 56448 49700 56500
rect 49752 56488 49758 56500
rect 50157 56491 50215 56497
rect 50157 56488 50169 56491
rect 49752 56460 50169 56488
rect 49752 56448 49758 56460
rect 50157 56457 50169 56460
rect 50203 56457 50215 56491
rect 51442 56488 51448 56500
rect 51403 56460 51448 56488
rect 50157 56451 50215 56457
rect 51442 56448 51448 56460
rect 51500 56448 51506 56500
rect 52822 56488 52828 56500
rect 52783 56460 52828 56488
rect 52822 56448 52828 56460
rect 52880 56448 52886 56500
rect 53834 56488 53840 56500
rect 53795 56460 53840 56488
rect 53834 56448 53840 56460
rect 53892 56448 53898 56500
rect 39853 56423 39911 56429
rect 39853 56389 39865 56423
rect 39899 56420 39911 56423
rect 43901 56423 43959 56429
rect 43901 56420 43913 56423
rect 39899 56392 43913 56420
rect 39899 56389 39911 56392
rect 39853 56383 39911 56389
rect 43901 56389 43913 56392
rect 43947 56389 43959 56423
rect 43901 56383 43959 56389
rect 43990 56380 43996 56432
rect 44048 56420 44054 56432
rect 44048 56392 44404 56420
rect 44048 56380 44054 56392
rect 39761 56355 39819 56361
rect 39761 56321 39773 56355
rect 39807 56321 39819 56355
rect 39942 56352 39948 56364
rect 39855 56324 39948 56352
rect 39761 56315 39819 56321
rect 39942 56312 39948 56324
rect 40000 56312 40006 56364
rect 40126 56361 40132 56364
rect 40083 56355 40132 56361
rect 40083 56321 40095 56355
rect 40129 56321 40132 56355
rect 40083 56315 40132 56321
rect 40126 56312 40132 56315
rect 40184 56312 40190 56364
rect 41138 56352 41144 56364
rect 41099 56324 41144 56352
rect 41138 56312 41144 56324
rect 41196 56312 41202 56364
rect 41966 56312 41972 56364
rect 42024 56352 42030 56364
rect 42061 56355 42119 56361
rect 42061 56352 42073 56355
rect 42024 56324 42073 56352
rect 42024 56312 42030 56324
rect 42061 56321 42073 56324
rect 42107 56321 42119 56355
rect 42061 56315 42119 56321
rect 43257 56355 43315 56361
rect 43257 56321 43269 56355
rect 43303 56352 43315 56355
rect 44082 56352 44088 56364
rect 43303 56324 43944 56352
rect 44043 56324 44088 56352
rect 43303 56321 43315 56324
rect 43257 56315 43315 56321
rect 34388 56256 34652 56284
rect 34388 56244 34394 56256
rect 34698 56244 34704 56296
rect 34756 56284 34762 56296
rect 34977 56287 35035 56293
rect 34977 56284 34989 56287
rect 34756 56256 34989 56284
rect 34756 56244 34762 56256
rect 34977 56253 34989 56256
rect 35023 56284 35035 56287
rect 35710 56284 35716 56296
rect 35023 56256 35716 56284
rect 35023 56253 35035 56256
rect 34977 56247 35035 56253
rect 35710 56244 35716 56256
rect 35768 56244 35774 56296
rect 37461 56287 37519 56293
rect 37461 56253 37473 56287
rect 37507 56284 37519 56287
rect 38013 56287 38071 56293
rect 38013 56284 38025 56287
rect 37507 56256 38025 56284
rect 37507 56253 37519 56256
rect 37461 56247 37519 56253
rect 38013 56253 38025 56256
rect 38059 56253 38071 56287
rect 38013 56247 38071 56253
rect 38194 56244 38200 56296
rect 38252 56284 38258 56296
rect 38473 56287 38531 56293
rect 38473 56284 38485 56287
rect 38252 56256 38485 56284
rect 38252 56244 38258 56256
rect 38473 56253 38485 56256
rect 38519 56253 38531 56287
rect 38473 56247 38531 56253
rect 38746 56244 38752 56296
rect 38804 56284 38810 56296
rect 39960 56284 39988 56312
rect 40218 56284 40224 56296
rect 38804 56256 39988 56284
rect 40179 56256 40224 56284
rect 38804 56244 38810 56256
rect 40218 56244 40224 56256
rect 40276 56244 40282 56296
rect 41417 56287 41475 56293
rect 41417 56253 41429 56287
rect 41463 56284 41475 56287
rect 41506 56284 41512 56296
rect 41463 56256 41512 56284
rect 41463 56253 41475 56256
rect 41417 56247 41475 56253
rect 41506 56244 41512 56256
rect 41564 56284 41570 56296
rect 42337 56287 42395 56293
rect 41564 56256 42104 56284
rect 41564 56244 41570 56256
rect 42076 56228 42104 56256
rect 42337 56253 42349 56287
rect 42383 56253 42395 56287
rect 43346 56284 43352 56296
rect 43307 56256 43352 56284
rect 42337 56247 42395 56253
rect 33594 56176 33600 56228
rect 33652 56216 33658 56228
rect 33652 56188 36308 56216
rect 33652 56176 33658 56188
rect 34698 56148 34704 56160
rect 33520 56120 34704 56148
rect 34698 56108 34704 56120
rect 34756 56108 34762 56160
rect 36280 56148 36308 56188
rect 37366 56176 37372 56228
rect 37424 56216 37430 56228
rect 38102 56216 38108 56228
rect 37424 56188 38108 56216
rect 37424 56176 37430 56188
rect 38102 56176 38108 56188
rect 38160 56176 38166 56228
rect 41874 56216 41880 56228
rect 41835 56188 41880 56216
rect 41874 56176 41880 56188
rect 41932 56176 41938 56228
rect 42058 56176 42064 56228
rect 42116 56176 42122 56228
rect 38933 56151 38991 56157
rect 38933 56148 38945 56151
rect 36280 56120 38945 56148
rect 38933 56117 38945 56120
rect 38979 56117 38991 56151
rect 38933 56111 38991 56117
rect 40402 56108 40408 56160
rect 40460 56148 40466 56160
rect 40954 56148 40960 56160
rect 40460 56120 40960 56148
rect 40460 56108 40466 56120
rect 40954 56108 40960 56120
rect 41012 56148 41018 56160
rect 41325 56151 41383 56157
rect 41325 56148 41337 56151
rect 41012 56120 41337 56148
rect 41012 56108 41018 56120
rect 41325 56117 41337 56120
rect 41371 56117 41383 56151
rect 42242 56148 42248 56160
rect 42203 56120 42248 56148
rect 41325 56111 41383 56117
rect 42242 56108 42248 56120
rect 42300 56108 42306 56160
rect 42352 56148 42380 56247
rect 43346 56244 43352 56256
rect 43404 56244 43410 56296
rect 43916 56284 43944 56324
rect 44082 56312 44088 56324
rect 44140 56312 44146 56364
rect 44376 56361 44404 56392
rect 44361 56355 44419 56361
rect 44361 56321 44373 56355
rect 44407 56321 44419 56355
rect 44361 56315 44419 56321
rect 45002 56312 45008 56364
rect 45060 56352 45066 56364
rect 45127 56355 45185 56361
rect 45127 56352 45139 56355
rect 45060 56324 45139 56352
rect 45060 56312 45066 56324
rect 45127 56321 45139 56324
rect 45173 56321 45185 56355
rect 45127 56315 45185 56321
rect 45278 56312 45284 56364
rect 45336 56352 45342 56364
rect 45336 56324 45381 56352
rect 45336 56312 45342 56324
rect 46474 56312 46480 56364
rect 46532 56352 46538 56364
rect 47029 56355 47087 56361
rect 47029 56352 47041 56355
rect 46532 56324 47041 56352
rect 46532 56312 46538 56324
rect 47029 56321 47041 56324
rect 47075 56321 47087 56355
rect 47029 56315 47087 56321
rect 47394 56312 47400 56364
rect 47452 56352 47458 56364
rect 47673 56355 47731 56361
rect 47673 56352 47685 56355
rect 47452 56324 47685 56352
rect 47452 56312 47458 56324
rect 47673 56321 47685 56324
rect 47719 56321 47731 56355
rect 47673 56315 47731 56321
rect 48774 56312 48780 56364
rect 48832 56352 48838 56364
rect 48869 56355 48927 56361
rect 48869 56352 48881 56355
rect 48832 56324 48881 56352
rect 48832 56312 48838 56324
rect 48869 56321 48881 56324
rect 48915 56321 48927 56355
rect 48869 56315 48927 56321
rect 49234 56312 49240 56364
rect 49292 56352 49298 56364
rect 49513 56355 49571 56361
rect 49513 56352 49525 56355
rect 49292 56324 49525 56352
rect 49292 56312 49298 56324
rect 49513 56321 49525 56324
rect 49559 56321 49571 56355
rect 49513 56315 49571 56321
rect 44266 56284 44272 56296
rect 43916 56256 44272 56284
rect 44266 56244 44272 56256
rect 44324 56244 44330 56296
rect 44634 56244 44640 56296
rect 44692 56284 44698 56296
rect 46385 56287 46443 56293
rect 46385 56284 46397 56287
rect 44692 56256 46397 56284
rect 44692 56244 44698 56256
rect 46385 56253 46397 56256
rect 46431 56253 46443 56287
rect 46385 56247 46443 56253
rect 42794 56176 42800 56228
rect 42852 56216 42858 56228
rect 42889 56219 42947 56225
rect 42889 56216 42901 56219
rect 42852 56188 42901 56216
rect 42852 56176 42858 56188
rect 42889 56185 42901 56188
rect 42935 56185 42947 56219
rect 42889 56179 42947 56185
rect 43254 56176 43260 56228
rect 43312 56216 43318 56228
rect 45741 56219 45799 56225
rect 45741 56216 45753 56219
rect 43312 56188 45753 56216
rect 43312 56176 43318 56188
rect 45741 56185 45753 56188
rect 45787 56185 45799 56219
rect 45741 56179 45799 56185
rect 42702 56148 42708 56160
rect 42352 56120 42708 56148
rect 42702 56108 42708 56120
rect 42760 56148 42766 56160
rect 44358 56148 44364 56160
rect 42760 56120 44364 56148
rect 42760 56108 42766 56120
rect 44358 56108 44364 56120
rect 44416 56108 44422 56160
rect 44542 56108 44548 56160
rect 44600 56148 44606 56160
rect 45097 56151 45155 56157
rect 45097 56148 45109 56151
rect 44600 56120 45109 56148
rect 44600 56108 44606 56120
rect 45097 56117 45109 56120
rect 45143 56117 45155 56151
rect 45097 56111 45155 56117
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 23934 55944 23940 55956
rect 23895 55916 23940 55944
rect 23934 55904 23940 55916
rect 23992 55904 23998 55956
rect 24765 55947 24823 55953
rect 24765 55913 24777 55947
rect 24811 55944 24823 55947
rect 25130 55944 25136 55956
rect 24811 55916 25136 55944
rect 24811 55913 24823 55916
rect 24765 55907 24823 55913
rect 25130 55904 25136 55916
rect 25188 55904 25194 55956
rect 25774 55904 25780 55956
rect 25832 55944 25838 55956
rect 26053 55947 26111 55953
rect 26053 55944 26065 55947
rect 25832 55916 26065 55944
rect 25832 55904 25838 55916
rect 26053 55913 26065 55916
rect 26099 55913 26111 55947
rect 26053 55907 26111 55913
rect 27341 55947 27399 55953
rect 27341 55913 27353 55947
rect 27387 55944 27399 55947
rect 28258 55944 28264 55956
rect 27387 55916 28264 55944
rect 27387 55913 27399 55916
rect 27341 55907 27399 55913
rect 28258 55904 28264 55916
rect 28316 55904 28322 55956
rect 28994 55904 29000 55956
rect 29052 55944 29058 55956
rect 35069 55947 35127 55953
rect 35069 55944 35081 55947
rect 29052 55916 35081 55944
rect 29052 55904 29058 55916
rect 35069 55913 35081 55916
rect 35115 55913 35127 55947
rect 35069 55907 35127 55913
rect 35434 55904 35440 55956
rect 35492 55944 35498 55956
rect 37182 55944 37188 55956
rect 35492 55916 37188 55944
rect 35492 55904 35498 55916
rect 37182 55904 37188 55916
rect 37240 55904 37246 55956
rect 37369 55947 37427 55953
rect 37369 55913 37381 55947
rect 37415 55944 37427 55947
rect 37458 55944 37464 55956
rect 37415 55916 37464 55944
rect 37415 55913 37427 55916
rect 37369 55907 37427 55913
rect 37458 55904 37464 55916
rect 37516 55904 37522 55956
rect 37829 55947 37887 55953
rect 37829 55913 37841 55947
rect 37875 55944 37887 55947
rect 38010 55944 38016 55956
rect 37875 55916 38016 55944
rect 37875 55913 37887 55916
rect 37829 55907 37887 55913
rect 38010 55904 38016 55916
rect 38068 55904 38074 55956
rect 38286 55904 38292 55956
rect 38344 55944 38350 55956
rect 40954 55944 40960 55956
rect 38344 55916 40960 55944
rect 38344 55904 38350 55916
rect 40954 55904 40960 55916
rect 41012 55904 41018 55956
rect 41601 55947 41659 55953
rect 41601 55913 41613 55947
rect 41647 55913 41659 55947
rect 44266 55944 44272 55956
rect 44227 55916 44272 55944
rect 41601 55907 41659 55913
rect 25148 55808 25176 55904
rect 25409 55879 25467 55885
rect 25409 55845 25421 55879
rect 25455 55876 25467 55879
rect 26694 55876 26700 55888
rect 25455 55848 26700 55876
rect 25455 55845 25467 55848
rect 25409 55839 25467 55845
rect 26694 55836 26700 55848
rect 26752 55836 26758 55888
rect 27890 55836 27896 55888
rect 27948 55876 27954 55888
rect 28629 55879 28687 55885
rect 28629 55876 28641 55879
rect 27948 55848 28641 55876
rect 27948 55836 27954 55848
rect 28629 55845 28641 55848
rect 28675 55845 28687 55879
rect 28629 55839 28687 55845
rect 28718 55836 28724 55888
rect 28776 55876 28782 55888
rect 31021 55879 31079 55885
rect 31021 55876 31033 55879
rect 28776 55848 31033 55876
rect 28776 55836 28782 55848
rect 31021 55845 31033 55848
rect 31067 55845 31079 55879
rect 31570 55876 31576 55888
rect 31021 55839 31079 55845
rect 31128 55848 31576 55876
rect 27801 55811 27859 55817
rect 27801 55808 27813 55811
rect 25148 55780 25912 55808
rect 24578 55740 24584 55752
rect 24539 55712 24584 55740
rect 24578 55700 24584 55712
rect 24636 55700 24642 55752
rect 25884 55749 25912 55780
rect 27172 55780 27813 55808
rect 27172 55749 27200 55780
rect 27801 55777 27813 55780
rect 27847 55808 27859 55811
rect 28997 55811 29055 55817
rect 27847 55780 28948 55808
rect 27847 55777 27859 55780
rect 27801 55771 27859 55777
rect 28920 55752 28948 55780
rect 28997 55777 29009 55811
rect 29043 55808 29055 55811
rect 29270 55808 29276 55820
rect 29043 55780 29276 55808
rect 29043 55777 29055 55780
rect 28997 55771 29055 55777
rect 29270 55768 29276 55780
rect 29328 55808 29334 55820
rect 31128 55808 31156 55848
rect 31570 55836 31576 55848
rect 31628 55836 31634 55888
rect 33042 55876 33048 55888
rect 33003 55848 33048 55876
rect 33042 55836 33048 55848
rect 33100 55836 33106 55888
rect 33686 55876 33692 55888
rect 33244 55848 33692 55876
rect 29328 55780 31156 55808
rect 29328 55768 29334 55780
rect 31294 55768 31300 55820
rect 31352 55768 31358 55820
rect 31662 55808 31668 55820
rect 31623 55780 31668 55808
rect 31662 55768 31668 55780
rect 31720 55768 31726 55820
rect 31206 55753 31264 55759
rect 25869 55743 25927 55749
rect 25869 55709 25881 55743
rect 25915 55709 25927 55743
rect 25869 55703 25927 55709
rect 27065 55743 27123 55749
rect 27065 55709 27077 55743
rect 27111 55709 27123 55743
rect 27065 55703 27123 55709
rect 27157 55743 27215 55749
rect 27157 55709 27169 55743
rect 27203 55709 27215 55743
rect 28810 55740 28816 55752
rect 27157 55703 27215 55709
rect 27264 55712 28816 55740
rect 27080 55672 27108 55703
rect 27264 55672 27292 55712
rect 28810 55700 28816 55712
rect 28868 55700 28874 55752
rect 28902 55700 28908 55752
rect 28960 55740 28966 55752
rect 29089 55743 29147 55749
rect 28960 55712 29005 55740
rect 28960 55700 28966 55712
rect 29089 55709 29101 55743
rect 29135 55740 29147 55743
rect 29730 55740 29736 55752
rect 29135 55712 29736 55740
rect 29135 55709 29147 55712
rect 29089 55703 29147 55709
rect 29730 55700 29736 55712
rect 29788 55700 29794 55752
rect 30282 55700 30288 55752
rect 30340 55740 30346 55752
rect 31206 55750 31218 55753
rect 30469 55743 30527 55749
rect 30340 55712 30385 55740
rect 30340 55700 30346 55712
rect 30469 55709 30481 55743
rect 30515 55740 30527 55743
rect 31128 55740 31218 55750
rect 30515 55722 31218 55740
rect 30515 55712 31156 55722
rect 31206 55719 31218 55722
rect 31252 55719 31264 55753
rect 31206 55713 31264 55719
rect 31312 55740 31340 55768
rect 31389 55743 31447 55749
rect 31389 55740 31401 55743
rect 31312 55712 31401 55740
rect 30515 55709 30527 55712
rect 30469 55703 30527 55709
rect 31389 55709 31401 55712
rect 31435 55740 31447 55743
rect 31938 55740 31944 55752
rect 31435 55712 31944 55740
rect 31435 55709 31447 55712
rect 31389 55703 31447 55709
rect 31938 55700 31944 55712
rect 31996 55700 32002 55752
rect 32309 55743 32367 55749
rect 32309 55709 32321 55743
rect 32355 55740 32367 55743
rect 32398 55740 32404 55752
rect 32355 55712 32404 55740
rect 32355 55709 32367 55712
rect 32309 55703 32367 55709
rect 32398 55700 32404 55712
rect 32456 55700 32462 55752
rect 32582 55740 32588 55752
rect 32543 55712 32588 55740
rect 32582 55700 32588 55712
rect 32640 55700 32646 55752
rect 33244 55749 33272 55848
rect 33686 55836 33692 55848
rect 33744 55836 33750 55888
rect 34054 55836 34060 55888
rect 34112 55876 34118 55888
rect 36538 55876 36544 55888
rect 34112 55848 36544 55876
rect 34112 55836 34118 55848
rect 36538 55836 36544 55848
rect 36596 55836 36602 55888
rect 36906 55836 36912 55888
rect 36964 55876 36970 55888
rect 39761 55879 39819 55885
rect 39761 55876 39773 55879
rect 36964 55848 39773 55876
rect 36964 55836 36970 55848
rect 39761 55845 39773 55848
rect 39807 55845 39819 55879
rect 41322 55876 41328 55888
rect 39761 55839 39819 55845
rect 39868 55848 41328 55876
rect 35437 55811 35495 55817
rect 35437 55777 35449 55811
rect 35483 55808 35495 55811
rect 35526 55808 35532 55820
rect 35483 55780 35532 55808
rect 35483 55777 35495 55780
rect 35437 55771 35495 55777
rect 35526 55768 35532 55780
rect 35584 55768 35590 55820
rect 36078 55768 36084 55820
rect 36136 55808 36142 55820
rect 36357 55811 36415 55817
rect 36357 55808 36369 55811
rect 36136 55780 36369 55808
rect 36136 55768 36142 55780
rect 36357 55777 36369 55780
rect 36403 55777 36415 55811
rect 39666 55808 39672 55820
rect 36357 55771 36415 55777
rect 38028 55780 39672 55808
rect 33244 55743 33306 55749
rect 33244 55712 33260 55743
rect 33248 55709 33260 55712
rect 33294 55709 33306 55743
rect 33248 55703 33306 55709
rect 33505 55743 33563 55749
rect 33505 55709 33517 55743
rect 33551 55740 33563 55743
rect 33778 55740 33784 55752
rect 33551 55712 33784 55740
rect 33551 55709 33563 55712
rect 33505 55703 33563 55709
rect 27080 55644 27292 55672
rect 27341 55675 27399 55681
rect 27341 55641 27353 55675
rect 27387 55641 27399 55675
rect 27982 55672 27988 55684
rect 27943 55644 27988 55672
rect 27341 55635 27399 55641
rect 23477 55607 23535 55613
rect 23477 55573 23489 55607
rect 23523 55604 23535 55607
rect 24486 55604 24492 55616
rect 23523 55576 24492 55604
rect 23523 55573 23535 55576
rect 23477 55567 23535 55573
rect 24486 55564 24492 55576
rect 24544 55564 24550 55616
rect 27356 55604 27384 55635
rect 27982 55632 27988 55644
rect 28040 55632 28046 55684
rect 28169 55675 28227 55681
rect 28169 55641 28181 55675
rect 28215 55672 28227 55675
rect 28994 55672 29000 55684
rect 28215 55644 29000 55672
rect 28215 55641 28227 55644
rect 28169 55635 28227 55641
rect 28994 55632 29000 55644
rect 29052 55632 29058 55684
rect 30098 55672 30104 55684
rect 30059 55644 30104 55672
rect 30098 55632 30104 55644
rect 30156 55632 30162 55684
rect 31297 55675 31355 55681
rect 31297 55641 31309 55675
rect 31343 55641 31355 55675
rect 31297 55635 31355 55641
rect 31527 55675 31585 55681
rect 31527 55641 31539 55675
rect 31573 55672 31585 55675
rect 31846 55672 31852 55684
rect 31573 55644 31852 55672
rect 31573 55641 31585 55644
rect 31527 55635 31585 55641
rect 29270 55604 29276 55616
rect 27356 55576 29276 55604
rect 29270 55564 29276 55576
rect 29328 55564 29334 55616
rect 31312 55604 31340 55635
rect 31846 55632 31852 55644
rect 31904 55632 31910 55684
rect 32490 55672 32496 55684
rect 32403 55644 32496 55672
rect 32490 55632 32496 55644
rect 32548 55672 32554 55684
rect 33520 55672 33548 55703
rect 33778 55700 33784 55712
rect 33836 55740 33842 55752
rect 34330 55740 34336 55752
rect 33836 55712 34336 55740
rect 33836 55700 33842 55712
rect 34330 55700 34336 55712
rect 34388 55700 34394 55752
rect 34425 55743 34483 55749
rect 34425 55709 34437 55743
rect 34471 55740 34483 55743
rect 34698 55740 34704 55752
rect 34471 55712 34704 55740
rect 34471 55709 34483 55712
rect 34425 55703 34483 55709
rect 34698 55700 34704 55712
rect 34756 55700 34762 55752
rect 35267 55743 35325 55749
rect 35267 55709 35279 55743
rect 35313 55709 35325 55743
rect 35267 55703 35325 55709
rect 35268 55672 35296 55703
rect 36262 55700 36268 55752
rect 36320 55740 36326 55752
rect 36541 55743 36599 55749
rect 36541 55740 36553 55743
rect 36320 55712 36553 55740
rect 36320 55700 36326 55712
rect 36541 55709 36553 55712
rect 36587 55709 36599 55743
rect 36814 55740 36820 55752
rect 36775 55712 36820 55740
rect 36541 55703 36599 55709
rect 36814 55700 36820 55712
rect 36872 55700 36878 55752
rect 38028 55749 38056 55780
rect 39666 55768 39672 55780
rect 39724 55768 39730 55820
rect 38013 55743 38071 55749
rect 38013 55709 38025 55743
rect 38059 55709 38071 55743
rect 38013 55703 38071 55709
rect 38105 55743 38163 55749
rect 38105 55709 38117 55743
rect 38151 55709 38163 55743
rect 38105 55703 38163 55709
rect 35710 55672 35716 55684
rect 32548 55644 33548 55672
rect 33980 55644 35716 55672
rect 32548 55632 32554 55644
rect 32125 55607 32183 55613
rect 32125 55604 32137 55607
rect 31312 55576 32137 55604
rect 32125 55573 32137 55576
rect 32171 55573 32183 55607
rect 32125 55567 32183 55573
rect 32766 55564 32772 55616
rect 32824 55604 32830 55616
rect 33413 55607 33471 55613
rect 33413 55604 33425 55607
rect 32824 55576 33425 55604
rect 32824 55564 32830 55576
rect 33413 55573 33425 55576
rect 33459 55604 33471 55607
rect 33980 55604 34008 55644
rect 35710 55632 35716 55644
rect 35768 55672 35774 55684
rect 38120 55672 38148 55703
rect 38194 55700 38200 55752
rect 38252 55740 38258 55752
rect 38289 55743 38347 55749
rect 38289 55740 38301 55743
rect 38252 55712 38301 55740
rect 38252 55700 38258 55712
rect 38289 55709 38301 55712
rect 38335 55709 38347 55743
rect 38289 55703 38347 55709
rect 38381 55743 38439 55749
rect 38381 55709 38393 55743
rect 38427 55740 38439 55743
rect 38746 55740 38752 55752
rect 38427 55712 38752 55740
rect 38427 55709 38439 55712
rect 38381 55703 38439 55709
rect 38746 55700 38752 55712
rect 38804 55700 38810 55752
rect 39206 55740 39212 55752
rect 39119 55712 39212 55740
rect 38470 55672 38476 55684
rect 35768 55644 36860 55672
rect 38120 55644 38476 55672
rect 35768 55632 35774 55644
rect 33459 55576 34008 55604
rect 34057 55607 34115 55613
rect 33459 55573 33471 55576
rect 33413 55567 33471 55573
rect 34057 55573 34069 55607
rect 34103 55604 34115 55607
rect 34514 55604 34520 55616
rect 34103 55576 34520 55604
rect 34103 55573 34115 55576
rect 34057 55567 34115 55573
rect 34514 55564 34520 55576
rect 34572 55564 34578 55616
rect 34790 55564 34796 55616
rect 34848 55604 34854 55616
rect 36078 55604 36084 55616
rect 34848 55576 36084 55604
rect 34848 55564 34854 55576
rect 36078 55564 36084 55576
rect 36136 55564 36142 55616
rect 36722 55604 36728 55616
rect 36683 55576 36728 55604
rect 36722 55564 36728 55576
rect 36780 55564 36786 55616
rect 36832 55604 36860 55644
rect 38470 55632 38476 55644
rect 38528 55672 38534 55684
rect 39132 55681 39160 55712
rect 39206 55700 39212 55712
rect 39264 55740 39270 55752
rect 39868 55740 39896 55848
rect 41322 55836 41328 55848
rect 41380 55836 41386 55888
rect 41616 55876 41644 55907
rect 44266 55904 44272 55916
rect 44324 55904 44330 55956
rect 44726 55904 44732 55956
rect 44784 55944 44790 55956
rect 45005 55947 45063 55953
rect 45005 55944 45017 55947
rect 44784 55916 45017 55944
rect 44784 55904 44790 55916
rect 45005 55913 45017 55916
rect 45051 55913 45063 55947
rect 45005 55907 45063 55913
rect 45094 55904 45100 55956
rect 45152 55944 45158 55956
rect 45649 55947 45707 55953
rect 45649 55944 45661 55947
rect 45152 55916 45661 55944
rect 45152 55904 45158 55916
rect 45649 55913 45661 55916
rect 45695 55913 45707 55947
rect 47578 55944 47584 55956
rect 47539 55916 47584 55944
rect 45649 55907 45707 55913
rect 47578 55904 47584 55916
rect 47636 55904 47642 55956
rect 48314 55944 48320 55956
rect 48275 55916 48320 55944
rect 48314 55904 48320 55916
rect 48372 55904 48378 55956
rect 41524 55848 41644 55876
rect 41046 55808 41052 55820
rect 40604 55780 41052 55808
rect 40604 55749 40632 55780
rect 41046 55768 41052 55780
rect 41104 55808 41110 55820
rect 41524 55808 41552 55848
rect 43622 55836 43628 55888
rect 43680 55876 43686 55888
rect 43680 55848 43725 55876
rect 43680 55836 43686 55848
rect 42245 55811 42303 55817
rect 42245 55808 42257 55811
rect 41104 55780 41552 55808
rect 41616 55780 42257 55808
rect 41104 55768 41110 55780
rect 39264 55712 39896 55740
rect 40589 55743 40647 55749
rect 39264 55700 39270 55712
rect 40589 55709 40601 55743
rect 40635 55709 40647 55743
rect 40862 55740 40868 55752
rect 40823 55712 40868 55740
rect 40589 55703 40647 55709
rect 40862 55700 40868 55712
rect 40920 55700 40926 55752
rect 40954 55700 40960 55752
rect 41012 55740 41018 55752
rect 41616 55740 41644 55780
rect 42245 55777 42257 55780
rect 42291 55777 42303 55811
rect 42245 55771 42303 55777
rect 43254 55768 43260 55820
rect 43312 55808 43318 55820
rect 43533 55811 43591 55817
rect 43533 55808 43545 55811
rect 43312 55780 43545 55808
rect 43312 55768 43318 55780
rect 43533 55777 43545 55780
rect 43579 55777 43591 55811
rect 44082 55808 44088 55820
rect 43533 55771 43591 55777
rect 43640 55780 44088 55808
rect 41012 55712 41644 55740
rect 41785 55743 41843 55749
rect 41012 55700 41018 55712
rect 41785 55709 41797 55743
rect 41831 55740 41843 55743
rect 41966 55740 41972 55752
rect 41831 55712 41972 55740
rect 41831 55709 41843 55712
rect 41785 55703 41843 55709
rect 38933 55675 38991 55681
rect 38933 55672 38945 55675
rect 38528 55644 38945 55672
rect 38528 55632 38534 55644
rect 38933 55641 38945 55644
rect 38979 55641 38991 55675
rect 38933 55635 38991 55641
rect 39117 55675 39175 55681
rect 39117 55641 39129 55675
rect 39163 55641 39175 55675
rect 39298 55672 39304 55684
rect 39259 55644 39304 55672
rect 39117 55635 39175 55641
rect 39298 55632 39304 55644
rect 39356 55632 39362 55684
rect 40773 55675 40831 55681
rect 40773 55641 40785 55675
rect 40819 55672 40831 55675
rect 41800 55672 41828 55703
rect 41966 55700 41972 55712
rect 42024 55700 42030 55752
rect 43438 55740 43444 55752
rect 43351 55712 43444 55740
rect 43438 55700 43444 55712
rect 43496 55740 43502 55752
rect 43640 55740 43668 55780
rect 44082 55768 44088 55780
rect 44140 55768 44146 55820
rect 44358 55768 44364 55820
rect 44416 55808 44422 55820
rect 45278 55808 45284 55820
rect 44416 55780 45284 55808
rect 44416 55768 44422 55780
rect 45278 55768 45284 55780
rect 45336 55768 45342 55820
rect 43496 55712 43668 55740
rect 43496 55700 43502 55712
rect 43714 55700 43720 55752
rect 43772 55740 43778 55752
rect 44542 55740 44548 55752
rect 43772 55712 44548 55740
rect 43772 55700 43778 55712
rect 44542 55700 44548 55712
rect 44600 55700 44606 55752
rect 40819 55644 41828 55672
rect 43257 55675 43315 55681
rect 40819 55641 40831 55644
rect 40773 55635 40831 55641
rect 43257 55641 43269 55675
rect 43303 55672 43315 55675
rect 43346 55672 43352 55684
rect 43303 55644 43352 55672
rect 43303 55641 43315 55644
rect 43257 55635 43315 55641
rect 43346 55632 43352 55644
rect 43404 55672 43410 55684
rect 44269 55675 44327 55681
rect 44269 55672 44281 55675
rect 43404 55644 44281 55672
rect 43404 55632 43410 55644
rect 44269 55641 44281 55644
rect 44315 55641 44327 55675
rect 44450 55672 44456 55684
rect 44411 55644 44456 55672
rect 44269 55635 44327 55641
rect 44450 55632 44456 55644
rect 44508 55632 44514 55684
rect 39022 55604 39028 55616
rect 36832 55576 39028 55604
rect 39022 55564 39028 55576
rect 39080 55564 39086 55616
rect 39758 55564 39764 55616
rect 39816 55604 39822 55616
rect 40405 55607 40463 55613
rect 40405 55604 40417 55607
rect 39816 55576 40417 55604
rect 39816 55564 39822 55576
rect 40405 55573 40417 55576
rect 40451 55573 40463 55607
rect 40405 55567 40463 55573
rect 40954 55564 40960 55616
rect 41012 55604 41018 55616
rect 41325 55607 41383 55613
rect 41325 55604 41337 55607
rect 41012 55576 41337 55604
rect 41012 55564 41018 55576
rect 41325 55573 41337 55576
rect 41371 55573 41383 55607
rect 41325 55567 41383 55573
rect 41506 55564 41512 55616
rect 41564 55604 41570 55616
rect 46750 55604 46756 55616
rect 41564 55576 46756 55604
rect 41564 55564 41570 55576
rect 46750 55564 46756 55576
rect 46808 55604 46814 55616
rect 46937 55607 46995 55613
rect 46937 55604 46949 55607
rect 46808 55576 46949 55604
rect 46808 55564 46814 55576
rect 46937 55573 46949 55576
rect 46983 55573 46995 55607
rect 46937 55567 46995 55573
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 25038 55360 25044 55412
rect 25096 55400 25102 55412
rect 25317 55403 25375 55409
rect 25317 55400 25329 55403
rect 25096 55372 25329 55400
rect 25096 55360 25102 55372
rect 25317 55369 25329 55372
rect 25363 55369 25375 55403
rect 25958 55400 25964 55412
rect 25919 55372 25964 55400
rect 25317 55363 25375 55369
rect 25958 55360 25964 55372
rect 26016 55360 26022 55412
rect 26789 55403 26847 55409
rect 26789 55369 26801 55403
rect 26835 55400 26847 55403
rect 26970 55400 26976 55412
rect 26835 55372 26976 55400
rect 26835 55369 26847 55372
rect 26789 55363 26847 55369
rect 26970 55360 26976 55372
rect 27028 55360 27034 55412
rect 27246 55360 27252 55412
rect 27304 55400 27310 55412
rect 27433 55403 27491 55409
rect 27433 55400 27445 55403
rect 27304 55372 27445 55400
rect 27304 55360 27310 55372
rect 27433 55369 27445 55372
rect 27479 55369 27491 55403
rect 27433 55363 27491 55369
rect 28537 55403 28595 55409
rect 28537 55369 28549 55403
rect 28583 55400 28595 55403
rect 29086 55400 29092 55412
rect 28583 55372 29092 55400
rect 28583 55369 28595 55372
rect 28537 55363 28595 55369
rect 29086 55360 29092 55372
rect 29144 55360 29150 55412
rect 30469 55403 30527 55409
rect 30469 55369 30481 55403
rect 30515 55369 30527 55403
rect 30469 55363 30527 55369
rect 31297 55403 31355 55409
rect 31297 55369 31309 55403
rect 31343 55400 31355 55403
rect 31343 55372 31524 55400
rect 31343 55369 31355 55372
rect 31297 55363 31355 55369
rect 28077 55335 28135 55341
rect 28077 55301 28089 55335
rect 28123 55332 28135 55335
rect 29362 55332 29368 55344
rect 28123 55304 29368 55332
rect 28123 55301 28135 55304
rect 28077 55295 28135 55301
rect 29362 55292 29368 55304
rect 29420 55332 29426 55344
rect 30484 55332 30512 55363
rect 31386 55332 31392 55344
rect 29420 55304 29776 55332
rect 30484 55304 31392 55332
rect 29420 55292 29426 55304
rect 25498 55264 25504 55276
rect 25459 55236 25504 55264
rect 25498 55224 25504 55236
rect 25556 55224 25562 55276
rect 26142 55264 26148 55276
rect 26103 55236 26148 55264
rect 26142 55224 26148 55236
rect 26200 55224 26206 55276
rect 26602 55264 26608 55276
rect 26563 55236 26608 55264
rect 26602 55224 26608 55236
rect 26660 55224 26666 55276
rect 26970 55224 26976 55276
rect 27028 55264 27034 55276
rect 27249 55267 27307 55273
rect 27249 55264 27261 55267
rect 27028 55236 27261 55264
rect 27028 55224 27034 55236
rect 27249 55233 27261 55236
rect 27295 55233 27307 55267
rect 27249 55227 27307 55233
rect 29457 55267 29515 55273
rect 29457 55233 29469 55267
rect 29503 55233 29515 55267
rect 29457 55227 29515 55233
rect 28810 55156 28816 55208
rect 28868 55196 28874 55208
rect 29273 55199 29331 55205
rect 29273 55196 29285 55199
rect 28868 55168 29285 55196
rect 28868 55156 28874 55168
rect 29273 55165 29285 55168
rect 29319 55165 29331 55199
rect 29472 55196 29500 55227
rect 29546 55224 29552 55276
rect 29604 55264 29610 55276
rect 29748 55273 29776 55304
rect 31386 55292 31392 55304
rect 31444 55292 31450 55344
rect 31496 55332 31524 55372
rect 31570 55360 31576 55412
rect 31628 55400 31634 55412
rect 35535 55403 35593 55409
rect 35535 55400 35547 55403
rect 31628 55372 35547 55400
rect 31628 55360 31634 55372
rect 35535 55369 35547 55372
rect 35581 55369 35593 55403
rect 35535 55363 35593 55369
rect 35621 55403 35679 55409
rect 35621 55369 35633 55403
rect 35667 55400 35679 55403
rect 35710 55400 35716 55412
rect 35667 55372 35716 55400
rect 35667 55369 35679 55372
rect 35621 55363 35679 55369
rect 35710 55360 35716 55372
rect 35768 55360 35774 55412
rect 35802 55360 35808 55412
rect 35860 55400 35866 55412
rect 37283 55403 37341 55409
rect 37283 55400 37295 55403
rect 35860 55372 37295 55400
rect 35860 55360 35866 55372
rect 37283 55369 37295 55372
rect 37329 55369 37341 55403
rect 37918 55400 37924 55412
rect 37879 55372 37924 55400
rect 37283 55363 37341 55369
rect 37918 55360 37924 55372
rect 37976 55360 37982 55412
rect 38289 55403 38347 55409
rect 38289 55369 38301 55403
rect 38335 55400 38347 55403
rect 38470 55400 38476 55412
rect 38335 55372 38476 55400
rect 38335 55369 38347 55372
rect 38289 55363 38347 55369
rect 38470 55360 38476 55372
rect 38528 55360 38534 55412
rect 39945 55403 40003 55409
rect 39945 55369 39957 55403
rect 39991 55400 40003 55403
rect 40862 55400 40868 55412
rect 39991 55372 40868 55400
rect 39991 55369 40003 55372
rect 39945 55363 40003 55369
rect 40862 55360 40868 55372
rect 40920 55360 40926 55412
rect 41125 55403 41183 55409
rect 41125 55369 41137 55403
rect 41171 55400 41183 55403
rect 41782 55400 41788 55412
rect 41171 55372 41788 55400
rect 41171 55369 41183 55372
rect 41125 55363 41183 55369
rect 41782 55360 41788 55372
rect 41840 55360 41846 55412
rect 43162 55400 43168 55412
rect 41892 55372 43168 55400
rect 31846 55332 31852 55344
rect 31496 55304 31852 55332
rect 31846 55292 31852 55304
rect 31904 55292 31910 55344
rect 34238 55292 34244 55344
rect 34296 55332 34302 55344
rect 34977 55335 35035 55341
rect 34296 55304 34836 55332
rect 34296 55292 34302 55304
rect 29733 55267 29791 55273
rect 29604 55236 29649 55264
rect 29604 55224 29610 55236
rect 29733 55233 29745 55267
rect 29779 55233 29791 55267
rect 29733 55227 29791 55233
rect 29825 55267 29883 55273
rect 29825 55233 29837 55267
rect 29871 55264 29883 55267
rect 30006 55264 30012 55276
rect 29871 55236 30012 55264
rect 29871 55233 29883 55236
rect 29825 55227 29883 55233
rect 30006 55224 30012 55236
rect 30064 55224 30070 55276
rect 30285 55267 30343 55273
rect 30285 55233 30297 55267
rect 30331 55264 30343 55267
rect 30466 55264 30472 55276
rect 30331 55236 30472 55264
rect 30331 55233 30343 55236
rect 30285 55227 30343 55233
rect 30466 55224 30472 55236
rect 30524 55224 30530 55276
rect 30926 55264 30932 55276
rect 30887 55236 30932 55264
rect 30926 55224 30932 55236
rect 30984 55224 30990 55276
rect 31110 55264 31116 55276
rect 31071 55236 31116 55264
rect 31110 55224 31116 55236
rect 31168 55224 31174 55276
rect 31754 55224 31760 55276
rect 31812 55264 31818 55276
rect 31941 55267 31999 55273
rect 31941 55264 31953 55267
rect 31812 55236 31953 55264
rect 31812 55224 31818 55236
rect 31941 55233 31953 55236
rect 31987 55233 31999 55267
rect 31941 55227 31999 55233
rect 32766 55224 32772 55276
rect 32824 55264 32830 55276
rect 33505 55267 33563 55273
rect 33505 55264 33517 55267
rect 32824 55236 33517 55264
rect 32824 55224 32830 55236
rect 33505 55233 33517 55236
rect 33551 55233 33563 55267
rect 34514 55264 34520 55276
rect 34475 55236 34520 55264
rect 33505 55227 33563 55233
rect 34514 55224 34520 55236
rect 34572 55224 34578 55276
rect 34808 55273 34836 55304
rect 34977 55301 34989 55335
rect 35023 55332 35035 55335
rect 35434 55332 35440 55344
rect 35023 55304 35440 55332
rect 35023 55301 35035 55304
rect 34977 55295 35035 55301
rect 35434 55292 35440 55304
rect 35492 55292 35498 55344
rect 37185 55335 37243 55341
rect 35544 55304 35848 55332
rect 34793 55267 34851 55273
rect 34793 55233 34805 55267
rect 34839 55264 34851 55267
rect 35544 55264 35572 55304
rect 34839 55236 35572 55264
rect 35713 55267 35771 55273
rect 34839 55233 34851 55236
rect 34793 55227 34851 55233
rect 35713 55233 35725 55267
rect 35759 55233 35771 55267
rect 35820 55264 35848 55304
rect 37185 55301 37197 55335
rect 37231 55332 37243 55335
rect 37550 55332 37556 55344
rect 37231 55304 37556 55332
rect 37231 55301 37243 55304
rect 37185 55295 37243 55301
rect 37550 55292 37556 55304
rect 37608 55292 37614 55344
rect 38746 55332 38752 55344
rect 38120 55304 38752 55332
rect 37366 55264 37372 55276
rect 35820 55236 37228 55264
rect 37327 55236 37372 55264
rect 35713 55227 35771 55233
rect 30944 55196 30972 55224
rect 29472 55168 30972 55196
rect 29273 55159 29331 55165
rect 32398 55156 32404 55208
rect 32456 55196 32462 55208
rect 34238 55196 34244 55208
rect 32456 55168 34244 55196
rect 32456 55156 32462 55168
rect 34238 55156 34244 55168
rect 34296 55156 34302 55208
rect 34532 55196 34560 55224
rect 35728 55196 35756 55227
rect 34532 55168 35756 55196
rect 35986 55156 35992 55208
rect 36044 55196 36050 55208
rect 36173 55199 36231 55205
rect 36173 55196 36185 55199
rect 36044 55168 36185 55196
rect 36044 55156 36050 55168
rect 36173 55165 36185 55168
rect 36219 55165 36231 55199
rect 37200 55196 37228 55236
rect 37366 55224 37372 55236
rect 37424 55224 37430 55276
rect 37461 55267 37519 55273
rect 37461 55233 37473 55267
rect 37507 55264 37519 55267
rect 38010 55264 38016 55276
rect 37507 55236 38016 55264
rect 37507 55233 37519 55236
rect 37461 55227 37519 55233
rect 38010 55224 38016 55236
rect 38068 55224 38074 55276
rect 38120 55273 38148 55304
rect 38746 55292 38752 55304
rect 38804 55332 38810 55344
rect 38930 55332 38936 55344
rect 38804 55304 38936 55332
rect 38804 55292 38810 55304
rect 38930 55292 38936 55304
rect 38988 55292 38994 55344
rect 41325 55335 41383 55341
rect 41325 55301 41337 55335
rect 41371 55332 41383 55335
rect 41892 55332 41920 55372
rect 43162 55360 43168 55372
rect 43220 55360 43226 55412
rect 45278 55360 45284 55412
rect 45336 55400 45342 55412
rect 46201 55403 46259 55409
rect 46201 55400 46213 55403
rect 45336 55372 46213 55400
rect 45336 55360 45342 55372
rect 46201 55369 46213 55372
rect 46247 55400 46259 55403
rect 54202 55400 54208 55412
rect 46247 55372 54208 55400
rect 46247 55369 46259 55372
rect 46201 55363 46259 55369
rect 54202 55360 54208 55372
rect 54260 55360 54266 55412
rect 43714 55332 43720 55344
rect 41371 55304 41920 55332
rect 42352 55304 43720 55332
rect 41371 55301 41383 55304
rect 41325 55295 41383 55301
rect 38105 55267 38163 55273
rect 38105 55233 38117 55267
rect 38151 55233 38163 55267
rect 38105 55227 38163 55233
rect 38381 55267 38439 55273
rect 38381 55233 38393 55267
rect 38427 55264 38439 55267
rect 39025 55267 39083 55273
rect 38427 55236 38792 55264
rect 38427 55233 38439 55236
rect 38381 55227 38439 55233
rect 38764 55208 38792 55236
rect 39025 55233 39037 55267
rect 39071 55264 39083 55267
rect 39206 55264 39212 55276
rect 39071 55236 39212 55264
rect 39071 55233 39083 55236
rect 39025 55227 39083 55233
rect 39206 55224 39212 55236
rect 39264 55224 39270 55276
rect 39574 55224 39580 55276
rect 39632 55264 39638 55276
rect 40034 55264 40040 55276
rect 39632 55236 40040 55264
rect 39632 55224 39638 55236
rect 40034 55224 40040 55236
rect 40092 55224 40098 55276
rect 40405 55267 40463 55273
rect 40405 55233 40417 55267
rect 40451 55264 40463 55267
rect 42058 55264 42064 55276
rect 40451 55236 42064 55264
rect 40451 55233 40463 55236
rect 40405 55227 40463 55233
rect 42058 55224 42064 55236
rect 42116 55224 42122 55276
rect 37274 55196 37280 55208
rect 37200 55168 37280 55196
rect 36173 55159 36231 55165
rect 37274 55156 37280 55168
rect 37332 55156 37338 55208
rect 38746 55156 38752 55208
rect 38804 55156 38810 55208
rect 38933 55199 38991 55205
rect 38933 55165 38945 55199
rect 38979 55165 38991 55199
rect 38933 55159 38991 55165
rect 28445 55131 28503 55137
rect 28445 55097 28457 55131
rect 28491 55128 28503 55131
rect 28902 55128 28908 55140
rect 28491 55100 28908 55128
rect 28491 55097 28503 55100
rect 28445 55091 28503 55097
rect 28902 55088 28908 55100
rect 28960 55088 28966 55140
rect 31294 55088 31300 55140
rect 31352 55128 31358 55140
rect 32582 55128 32588 55140
rect 31352 55100 32588 55128
rect 31352 55088 31358 55100
rect 32582 55088 32588 55100
rect 32640 55088 32646 55140
rect 34422 55088 34428 55140
rect 34480 55128 34486 55140
rect 34609 55131 34667 55137
rect 34609 55128 34621 55131
rect 34480 55100 34621 55128
rect 34480 55088 34486 55100
rect 34609 55097 34621 55100
rect 34655 55097 34667 55131
rect 34609 55091 34667 55097
rect 34698 55088 34704 55140
rect 34756 55128 34762 55140
rect 38948 55128 38976 55159
rect 41690 55156 41696 55208
rect 41748 55196 41754 55208
rect 41969 55199 42027 55205
rect 41969 55196 41981 55199
rect 41748 55168 41981 55196
rect 41748 55156 41754 55168
rect 41969 55165 41981 55168
rect 42015 55196 42027 55199
rect 42352 55196 42380 55304
rect 43714 55292 43720 55304
rect 43772 55332 43778 55344
rect 43772 55304 44128 55332
rect 43772 55292 43778 55304
rect 43257 55267 43315 55273
rect 43257 55233 43269 55267
rect 43303 55264 43315 55267
rect 43438 55264 43444 55276
rect 43303 55236 43444 55264
rect 43303 55233 43315 55236
rect 43257 55227 43315 55233
rect 43438 55224 43444 55236
rect 43496 55224 43502 55276
rect 44100 55273 44128 55304
rect 44085 55267 44143 55273
rect 44085 55233 44097 55267
rect 44131 55233 44143 55267
rect 44085 55227 44143 55233
rect 44174 55224 44180 55276
rect 44232 55264 44238 55276
rect 45097 55267 45155 55273
rect 45097 55264 45109 55267
rect 44232 55236 45109 55264
rect 44232 55224 44238 55236
rect 45097 55233 45109 55236
rect 45143 55264 45155 55267
rect 45557 55267 45615 55273
rect 45557 55264 45569 55267
rect 45143 55236 45569 55264
rect 45143 55233 45155 55236
rect 45097 55227 45155 55233
rect 45557 55233 45569 55236
rect 45603 55233 45615 55267
rect 45557 55227 45615 55233
rect 42015 55168 42380 55196
rect 42015 55165 42027 55168
rect 41969 55159 42027 55165
rect 42426 55156 42432 55208
rect 42484 55196 42490 55208
rect 43349 55199 43407 55205
rect 42484 55168 43300 55196
rect 42484 55156 42490 55168
rect 39114 55128 39120 55140
rect 34756 55100 34849 55128
rect 38948 55100 39120 55128
rect 34756 55088 34762 55100
rect 39114 55088 39120 55100
rect 39172 55128 39178 55140
rect 39298 55128 39304 55140
rect 39172 55100 39304 55128
rect 39172 55088 39178 55100
rect 39298 55088 39304 55100
rect 39356 55128 39362 55140
rect 42889 55131 42947 55137
rect 42889 55128 42901 55131
rect 39356 55100 42901 55128
rect 39356 55088 39362 55100
rect 42889 55097 42901 55100
rect 42935 55097 42947 55131
rect 43272 55128 43300 55168
rect 43349 55165 43361 55199
rect 43395 55196 43407 55199
rect 43901 55199 43959 55205
rect 43901 55196 43913 55199
rect 43395 55168 43913 55196
rect 43395 55165 43407 55168
rect 43349 55159 43407 55165
rect 43901 55165 43913 55168
rect 43947 55165 43959 55199
rect 43901 55159 43959 55165
rect 44361 55199 44419 55205
rect 44361 55165 44373 55199
rect 44407 55196 44419 55199
rect 45922 55196 45928 55208
rect 44407 55168 45928 55196
rect 44407 55165 44419 55168
rect 44361 55159 44419 55165
rect 43622 55128 43628 55140
rect 43272 55100 43628 55128
rect 42889 55091 42947 55097
rect 43622 55088 43628 55100
rect 43680 55128 43686 55140
rect 44269 55131 44327 55137
rect 44269 55128 44281 55131
rect 43680 55100 44281 55128
rect 43680 55088 43686 55100
rect 44269 55097 44281 55100
rect 44315 55097 44327 55131
rect 44269 55091 44327 55097
rect 24029 55063 24087 55069
rect 24029 55029 24041 55063
rect 24075 55060 24087 55063
rect 24578 55060 24584 55072
rect 24075 55032 24584 55060
rect 24075 55029 24087 55032
rect 24029 55023 24087 55029
rect 24578 55020 24584 55032
rect 24636 55020 24642 55072
rect 32030 55060 32036 55072
rect 31991 55032 32036 55060
rect 32030 55020 32036 55032
rect 32088 55020 32094 55072
rect 32398 55060 32404 55072
rect 32359 55032 32404 55060
rect 32398 55020 32404 55032
rect 32456 55020 32462 55072
rect 33042 55060 33048 55072
rect 33003 55032 33048 55060
rect 33042 55020 33048 55032
rect 33100 55020 33106 55072
rect 33413 55063 33471 55069
rect 33413 55029 33425 55063
rect 33459 55060 33471 55063
rect 33594 55060 33600 55072
rect 33459 55032 33600 55060
rect 33459 55029 33471 55032
rect 33413 55023 33471 55029
rect 33594 55020 33600 55032
rect 33652 55020 33658 55072
rect 33962 55020 33968 55072
rect 34020 55060 34026 55072
rect 34716 55060 34744 55088
rect 34020 55032 34744 55060
rect 39393 55063 39451 55069
rect 34020 55020 34026 55032
rect 39393 55029 39405 55063
rect 39439 55060 39451 55063
rect 39574 55060 39580 55072
rect 39439 55032 39580 55060
rect 39439 55029 39451 55032
rect 39393 55023 39451 55029
rect 39574 55020 39580 55032
rect 39632 55020 39638 55072
rect 40313 55063 40371 55069
rect 40313 55029 40325 55063
rect 40359 55060 40371 55063
rect 40402 55060 40408 55072
rect 40359 55032 40408 55060
rect 40359 55029 40371 55032
rect 40313 55023 40371 55029
rect 40402 55020 40408 55032
rect 40460 55020 40466 55072
rect 40957 55063 41015 55069
rect 40957 55029 40969 55063
rect 41003 55060 41015 55063
rect 41046 55060 41052 55072
rect 41003 55032 41052 55060
rect 41003 55029 41015 55032
rect 40957 55023 41015 55029
rect 41046 55020 41052 55032
rect 41104 55020 41110 55072
rect 41141 55063 41199 55069
rect 41141 55029 41153 55063
rect 41187 55060 41199 55063
rect 41874 55060 41880 55072
rect 41187 55032 41880 55060
rect 41187 55029 41199 55032
rect 41141 55023 41199 55029
rect 41874 55020 41880 55032
rect 41932 55020 41938 55072
rect 42058 55020 42064 55072
rect 42116 55060 42122 55072
rect 43254 55060 43260 55072
rect 42116 55032 43260 55060
rect 42116 55020 42122 55032
rect 43254 55020 43260 55032
rect 43312 55060 43318 55072
rect 44376 55060 44404 55159
rect 45922 55156 45928 55168
rect 45980 55156 45986 55208
rect 44910 55060 44916 55072
rect 43312 55032 44404 55060
rect 44871 55032 44916 55060
rect 43312 55020 43318 55032
rect 44910 55020 44916 55032
rect 44968 55020 44974 55072
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 25314 54816 25320 54868
rect 25372 54856 25378 54868
rect 25409 54859 25467 54865
rect 25409 54856 25421 54859
rect 25372 54828 25421 54856
rect 25372 54816 25378 54828
rect 25409 54825 25421 54828
rect 25455 54825 25467 54859
rect 25409 54819 25467 54825
rect 27709 54859 27767 54865
rect 27709 54825 27721 54859
rect 27755 54856 27767 54859
rect 28074 54856 28080 54868
rect 27755 54828 28080 54856
rect 27755 54825 27767 54828
rect 27709 54819 27767 54825
rect 28074 54816 28080 54828
rect 28132 54816 28138 54868
rect 28350 54856 28356 54868
rect 28311 54828 28356 54856
rect 28350 54816 28356 54828
rect 28408 54816 28414 54868
rect 30466 54816 30472 54868
rect 30524 54816 30530 54868
rect 31021 54859 31079 54865
rect 31021 54825 31033 54859
rect 31067 54856 31079 54859
rect 31110 54856 31116 54868
rect 31067 54828 31116 54856
rect 31067 54825 31079 54828
rect 31021 54819 31079 54825
rect 31110 54816 31116 54828
rect 31168 54816 31174 54868
rect 33137 54859 33195 54865
rect 33137 54856 33149 54859
rect 31220 54828 33149 54856
rect 29270 54748 29276 54800
rect 29328 54788 29334 54800
rect 29365 54791 29423 54797
rect 29365 54788 29377 54791
rect 29328 54760 29377 54788
rect 29328 54748 29334 54760
rect 29365 54757 29377 54760
rect 29411 54788 29423 54791
rect 29638 54788 29644 54800
rect 29411 54760 29644 54788
rect 29411 54757 29423 54760
rect 29365 54751 29423 54757
rect 29638 54748 29644 54760
rect 29696 54748 29702 54800
rect 30484 54788 30512 54816
rect 31220 54788 31248 54828
rect 33137 54825 33149 54828
rect 33183 54825 33195 54859
rect 33137 54819 33195 54825
rect 33318 54816 33324 54868
rect 33376 54856 33382 54868
rect 35897 54859 35955 54865
rect 35897 54856 35909 54859
rect 33376 54828 35909 54856
rect 33376 54816 33382 54828
rect 35897 54825 35909 54828
rect 35943 54825 35955 54859
rect 36538 54856 36544 54868
rect 36499 54828 36544 54856
rect 35897 54819 35955 54825
rect 36538 54816 36544 54828
rect 36596 54816 36602 54868
rect 37182 54856 37188 54868
rect 37143 54828 37188 54856
rect 37182 54816 37188 54828
rect 37240 54816 37246 54868
rect 38013 54859 38071 54865
rect 38013 54825 38025 54859
rect 38059 54856 38071 54859
rect 38194 54856 38200 54868
rect 38059 54828 38200 54856
rect 38059 54825 38071 54828
rect 38013 54819 38071 54825
rect 38194 54816 38200 54828
rect 38252 54816 38258 54868
rect 38930 54856 38936 54868
rect 38891 54828 38936 54856
rect 38930 54816 38936 54828
rect 38988 54816 38994 54868
rect 40126 54856 40132 54868
rect 40087 54828 40132 54856
rect 40126 54816 40132 54828
rect 40184 54816 40190 54868
rect 41966 54816 41972 54868
rect 42024 54856 42030 54868
rect 42245 54859 42303 54865
rect 42245 54856 42257 54859
rect 42024 54828 42257 54856
rect 42024 54816 42030 54828
rect 42245 54825 42257 54828
rect 42291 54825 42303 54859
rect 42886 54856 42892 54868
rect 42847 54828 42892 54856
rect 42245 54819 42303 54825
rect 42886 54816 42892 54828
rect 42944 54816 42950 54868
rect 43530 54856 43536 54868
rect 43491 54828 43536 54856
rect 43530 54816 43536 54828
rect 43588 54816 43594 54868
rect 30484 54760 31248 54788
rect 31754 54748 31760 54800
rect 31812 54788 31818 54800
rect 32677 54791 32735 54797
rect 31812 54760 32536 54788
rect 31812 54748 31818 54760
rect 28626 54720 28632 54732
rect 28184 54692 28632 54720
rect 28184 54661 28212 54692
rect 28626 54680 28632 54692
rect 28684 54680 28690 54732
rect 29086 54720 29092 54732
rect 29047 54692 29092 54720
rect 29086 54680 29092 54692
rect 29144 54680 29150 54732
rect 30098 54680 30104 54732
rect 30156 54720 30162 54732
rect 31481 54723 31539 54729
rect 30156 54692 30512 54720
rect 30156 54680 30162 54692
rect 28169 54655 28227 54661
rect 28169 54621 28181 54655
rect 28215 54621 28227 54655
rect 28169 54615 28227 54621
rect 28353 54655 28411 54661
rect 28353 54621 28365 54655
rect 28399 54652 28411 54655
rect 28534 54652 28540 54664
rect 28399 54624 28540 54652
rect 28399 54621 28411 54624
rect 28353 54615 28411 54621
rect 28534 54612 28540 54624
rect 28592 54612 28598 54664
rect 28997 54655 29055 54661
rect 28997 54621 29009 54655
rect 29043 54652 29055 54655
rect 29362 54652 29368 54664
rect 29043 54624 29368 54652
rect 29043 54621 29055 54624
rect 28997 54615 29055 54621
rect 29362 54612 29368 54624
rect 29420 54612 29426 54664
rect 30484 54661 30512 54692
rect 31481 54689 31493 54723
rect 31527 54689 31539 54723
rect 32398 54720 32404 54732
rect 32359 54692 32404 54720
rect 31481 54683 31539 54689
rect 30285 54655 30343 54661
rect 30285 54621 30297 54655
rect 30331 54621 30343 54655
rect 30285 54615 30343 54621
rect 30469 54655 30527 54661
rect 30469 54621 30481 54655
rect 30515 54652 30527 54655
rect 31294 54652 31300 54664
rect 30515 54624 31300 54652
rect 30515 54621 30527 54624
rect 30469 54615 30527 54621
rect 30300 54584 30328 54615
rect 31294 54612 31300 54624
rect 31352 54652 31358 54664
rect 31389 54655 31447 54661
rect 31389 54652 31401 54655
rect 31352 54624 31401 54652
rect 31352 54612 31358 54624
rect 31389 54621 31401 54624
rect 31435 54621 31447 54655
rect 31389 54615 31447 54621
rect 31496 54584 31524 54683
rect 32398 54680 32404 54692
rect 32456 54680 32462 54732
rect 32508 54720 32536 54760
rect 32677 54757 32689 54791
rect 32723 54788 32735 54791
rect 33410 54788 33416 54800
rect 32723 54760 33416 54788
rect 32723 54757 32735 54760
rect 32677 54751 32735 54757
rect 33410 54748 33416 54760
rect 33468 54748 33474 54800
rect 38562 54788 38568 54800
rect 38212 54760 38568 54788
rect 33873 54723 33931 54729
rect 32508 54692 33824 54720
rect 32309 54655 32367 54661
rect 32309 54621 32321 54655
rect 32355 54652 32367 54655
rect 33042 54652 33048 54664
rect 32355 54624 33048 54652
rect 32355 54621 32367 54624
rect 32309 54615 32367 54621
rect 33042 54612 33048 54624
rect 33100 54612 33106 54664
rect 33796 54652 33824 54692
rect 33873 54689 33885 54723
rect 33919 54720 33931 54723
rect 34514 54720 34520 54732
rect 33919 54692 34520 54720
rect 33919 54689 33931 54692
rect 33873 54683 33931 54689
rect 34514 54680 34520 54692
rect 34572 54680 34578 54732
rect 34606 54680 34612 54732
rect 34664 54720 34670 54732
rect 34974 54720 34980 54732
rect 34664 54692 34980 54720
rect 34664 54680 34670 54692
rect 34974 54680 34980 54692
rect 35032 54720 35038 54732
rect 35032 54692 35296 54720
rect 35032 54680 35038 54692
rect 33962 54652 33968 54664
rect 33796 54624 33968 54652
rect 33962 54612 33968 54624
rect 34020 54612 34026 54664
rect 34333 54655 34391 54661
rect 34333 54621 34345 54655
rect 34379 54652 34391 54655
rect 34422 54652 34428 54664
rect 34379 54624 34428 54652
rect 34379 54621 34391 54624
rect 34333 54615 34391 54621
rect 34422 54612 34428 54624
rect 34480 54612 34486 54664
rect 34532 54652 34560 54680
rect 34698 54652 34704 54664
rect 34532 54624 34704 54652
rect 34698 54612 34704 54624
rect 34756 54652 34762 54664
rect 35268 54661 35296 54692
rect 35161 54655 35219 54661
rect 35161 54652 35173 54655
rect 34756 54624 35173 54652
rect 34756 54612 34762 54624
rect 35161 54621 35173 54624
rect 35207 54621 35219 54655
rect 35161 54615 35219 54621
rect 35253 54655 35311 54661
rect 35253 54621 35265 54655
rect 35299 54621 35311 54655
rect 35253 54615 35311 54621
rect 35345 54655 35403 54661
rect 35345 54621 35357 54655
rect 35391 54621 35403 54655
rect 35345 54615 35403 54621
rect 33502 54584 33508 54596
rect 30300 54556 33508 54584
rect 30484 54528 30512 54556
rect 33502 54544 33508 54556
rect 33560 54544 33566 54596
rect 34440 54584 34468 54612
rect 34882 54584 34888 54596
rect 34440 54556 34888 54584
rect 34882 54544 34888 54556
rect 34940 54584 34946 54596
rect 35360 54584 35388 54615
rect 35894 54612 35900 54664
rect 35952 54652 35958 54664
rect 38212 54661 38240 54760
rect 38562 54748 38568 54760
rect 38620 54788 38626 54800
rect 42794 54788 42800 54800
rect 38620 54760 42800 54788
rect 38620 54748 38626 54760
rect 42794 54748 42800 54760
rect 42852 54748 42858 54800
rect 38378 54720 38384 54732
rect 38291 54692 38384 54720
rect 38378 54680 38384 54692
rect 38436 54720 38442 54732
rect 40862 54720 40868 54732
rect 38436 54692 40080 54720
rect 40823 54692 40868 54720
rect 38436 54680 38442 54692
rect 36081 54655 36139 54661
rect 36081 54652 36093 54655
rect 35952 54624 36093 54652
rect 35952 54612 35958 54624
rect 36081 54621 36093 54624
rect 36127 54621 36139 54655
rect 36081 54615 36139 54621
rect 38197 54655 38255 54661
rect 38197 54621 38209 54655
rect 38243 54621 38255 54655
rect 39114 54652 39120 54664
rect 39075 54624 39120 54652
rect 38197 54615 38255 54621
rect 39114 54612 39120 54624
rect 39172 54612 39178 54664
rect 39206 54612 39212 54664
rect 39264 54652 39270 54664
rect 39264 54624 39309 54652
rect 39264 54612 39270 54624
rect 39574 54612 39580 54664
rect 39632 54652 39638 54664
rect 39945 54655 40003 54661
rect 39945 54652 39957 54655
rect 39632 54624 39957 54652
rect 39632 54612 39638 54624
rect 39945 54621 39957 54624
rect 39991 54621 40003 54655
rect 39945 54615 40003 54621
rect 34940 54556 35388 54584
rect 34940 54544 34946 54556
rect 38746 54544 38752 54596
rect 38804 54584 38810 54596
rect 39758 54584 39764 54596
rect 38804 54556 39764 54584
rect 38804 54544 38810 54556
rect 39758 54544 39764 54556
rect 39816 54544 39822 54596
rect 40052 54584 40080 54692
rect 40862 54680 40868 54692
rect 40920 54680 40926 54732
rect 40954 54652 40960 54664
rect 40915 54624 40960 54652
rect 40954 54612 40960 54624
rect 41012 54612 41018 54664
rect 41782 54652 41788 54664
rect 41743 54624 41788 54652
rect 41782 54612 41788 54624
rect 41840 54612 41846 54664
rect 41874 54612 41880 54664
rect 41932 54652 41938 54664
rect 42061 54655 42119 54661
rect 41932 54624 41977 54652
rect 41932 54612 41938 54624
rect 42061 54621 42073 54655
rect 42107 54652 42119 54655
rect 43162 54652 43168 54664
rect 42107 54624 43168 54652
rect 42107 54621 42119 54624
rect 42061 54615 42119 54621
rect 43162 54612 43168 54624
rect 43220 54612 43226 54664
rect 44910 54584 44916 54596
rect 40052 54556 44916 54584
rect 44910 54544 44916 54556
rect 44968 54544 44974 54596
rect 24578 54516 24584 54528
rect 24491 54488 24584 54516
rect 24578 54476 24584 54488
rect 24636 54516 24642 54528
rect 26418 54516 26424 54528
rect 24636 54488 26424 54516
rect 24636 54476 24642 54488
rect 26418 54476 26424 54488
rect 26476 54476 26482 54528
rect 30006 54476 30012 54528
rect 30064 54516 30070 54528
rect 30101 54519 30159 54525
rect 30101 54516 30113 54519
rect 30064 54488 30113 54516
rect 30064 54476 30070 54488
rect 30101 54485 30113 54488
rect 30147 54485 30159 54519
rect 30101 54479 30159 54485
rect 30466 54476 30472 54528
rect 30524 54476 30530 54528
rect 33134 54476 33140 54528
rect 33192 54516 33198 54528
rect 33689 54519 33747 54525
rect 33689 54516 33701 54519
rect 33192 54488 33701 54516
rect 33192 54476 33198 54488
rect 33689 54485 33701 54488
rect 33735 54485 33747 54519
rect 33689 54479 33747 54485
rect 34422 54476 34428 54528
rect 34480 54516 34486 54528
rect 34977 54519 35035 54525
rect 34977 54516 34989 54519
rect 34480 54488 34989 54516
rect 34480 54476 34486 54488
rect 34977 54485 34989 54488
rect 35023 54485 35035 54519
rect 34977 54479 35035 54485
rect 41325 54519 41383 54525
rect 41325 54485 41337 54519
rect 41371 54516 41383 54519
rect 42242 54516 42248 54528
rect 41371 54488 42248 54516
rect 41371 54485 41383 54488
rect 41325 54479 41383 54485
rect 42242 54476 42248 54488
rect 42300 54476 42306 54528
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 25866 54312 25872 54324
rect 25827 54284 25872 54312
rect 25866 54272 25872 54284
rect 25924 54312 25930 54324
rect 26421 54315 26479 54321
rect 26421 54312 26433 54315
rect 25924 54284 26433 54312
rect 25924 54272 25930 54284
rect 26421 54281 26433 54284
rect 26467 54281 26479 54315
rect 26421 54275 26479 54281
rect 27341 54315 27399 54321
rect 27341 54281 27353 54315
rect 27387 54312 27399 54315
rect 27614 54312 27620 54324
rect 27387 54284 27620 54312
rect 27387 54281 27399 54284
rect 27341 54275 27399 54281
rect 27614 54272 27620 54284
rect 27672 54272 27678 54324
rect 29546 54312 29552 54324
rect 29507 54284 29552 54312
rect 29546 54272 29552 54284
rect 29604 54312 29610 54324
rect 30101 54315 30159 54321
rect 30101 54312 30113 54315
rect 29604 54284 30113 54312
rect 29604 54272 29610 54284
rect 30101 54281 30113 54284
rect 30147 54281 30159 54315
rect 30101 54275 30159 54281
rect 31021 54315 31079 54321
rect 31021 54281 31033 54315
rect 31067 54312 31079 54315
rect 31110 54312 31116 54324
rect 31067 54284 31116 54312
rect 31067 54281 31079 54284
rect 31021 54275 31079 54281
rect 31110 54272 31116 54284
rect 31168 54272 31174 54324
rect 32401 54315 32459 54321
rect 32401 54281 32413 54315
rect 32447 54312 32459 54315
rect 32766 54312 32772 54324
rect 32447 54284 32772 54312
rect 32447 54281 32459 54284
rect 32401 54275 32459 54281
rect 32766 54272 32772 54284
rect 32824 54272 32830 54324
rect 33502 54312 33508 54324
rect 33463 54284 33508 54312
rect 33502 54272 33508 54284
rect 33560 54272 33566 54324
rect 33686 54272 33692 54324
rect 33744 54312 33750 54324
rect 35529 54315 35587 54321
rect 35529 54312 35541 54315
rect 33744 54284 35541 54312
rect 33744 54272 33750 54284
rect 35529 54281 35541 54284
rect 35575 54281 35587 54315
rect 35529 54275 35587 54281
rect 37366 54272 37372 54324
rect 37424 54312 37430 54324
rect 38197 54315 38255 54321
rect 38197 54312 38209 54315
rect 37424 54284 38209 54312
rect 37424 54272 37430 54284
rect 38197 54281 38209 54284
rect 38243 54281 38255 54315
rect 39574 54312 39580 54324
rect 39535 54284 39580 54312
rect 38197 54275 38255 54281
rect 39574 54272 39580 54284
rect 39632 54272 39638 54324
rect 40402 54272 40408 54324
rect 40460 54312 40466 54324
rect 41141 54315 41199 54321
rect 41141 54312 41153 54315
rect 40460 54284 41153 54312
rect 40460 54272 40466 54284
rect 41141 54281 41153 54284
rect 41187 54281 41199 54315
rect 41141 54275 41199 54281
rect 41785 54315 41843 54321
rect 41785 54281 41797 54315
rect 41831 54312 41843 54315
rect 41874 54312 41880 54324
rect 41831 54284 41880 54312
rect 41831 54281 41843 54284
rect 41785 54275 41843 54281
rect 41874 54272 41880 54284
rect 41932 54272 41938 54324
rect 42058 54272 42064 54324
rect 42116 54272 42122 54324
rect 42702 54272 42708 54324
rect 42760 54312 42766 54324
rect 42797 54315 42855 54321
rect 42797 54312 42809 54315
rect 42760 54284 42809 54312
rect 42760 54272 42766 54284
rect 42797 54281 42809 54284
rect 42843 54281 42855 54315
rect 42797 54275 42855 54281
rect 29365 54247 29423 54253
rect 29365 54213 29377 54247
rect 29411 54244 29423 54247
rect 30006 54244 30012 54256
rect 29411 54216 30012 54244
rect 29411 54213 29423 54216
rect 29365 54207 29423 54213
rect 30006 54204 30012 54216
rect 30064 54204 30070 54256
rect 30466 54244 30472 54256
rect 30427 54216 30472 54244
rect 30466 54204 30472 54216
rect 30524 54204 30530 54256
rect 31205 54247 31263 54253
rect 31205 54213 31217 54247
rect 31251 54244 31263 54247
rect 31938 54244 31944 54256
rect 31251 54216 31944 54244
rect 31251 54213 31263 54216
rect 31205 54207 31263 54213
rect 31938 54204 31944 54216
rect 31996 54204 32002 54256
rect 33594 54244 33600 54256
rect 32232 54216 33600 54244
rect 27893 54179 27951 54185
rect 27893 54145 27905 54179
rect 27939 54176 27951 54179
rect 28353 54179 28411 54185
rect 28353 54176 28365 54179
rect 27939 54148 28365 54176
rect 27939 54145 27951 54148
rect 27893 54139 27951 54145
rect 28353 54145 28365 54148
rect 28399 54176 28411 54179
rect 28994 54176 29000 54188
rect 28399 54148 29000 54176
rect 28399 54145 28411 54148
rect 28353 54139 28411 54145
rect 28994 54136 29000 54148
rect 29052 54136 29058 54188
rect 29641 54179 29699 54185
rect 29641 54145 29653 54179
rect 29687 54145 29699 54179
rect 29641 54139 29699 54145
rect 29656 54108 29684 54139
rect 30098 54136 30104 54188
rect 30156 54176 30162 54188
rect 30285 54179 30343 54185
rect 30285 54176 30297 54179
rect 30156 54148 30297 54176
rect 30156 54136 30162 54148
rect 30285 54145 30297 54148
rect 30331 54145 30343 54179
rect 30926 54176 30932 54188
rect 30839 54148 30932 54176
rect 30285 54139 30343 54145
rect 30926 54136 30932 54148
rect 30984 54136 30990 54188
rect 32232 54185 32260 54216
rect 33594 54204 33600 54216
rect 33652 54204 33658 54256
rect 37458 54204 37464 54256
rect 37516 54244 37522 54256
rect 37645 54247 37703 54253
rect 37645 54244 37657 54247
rect 37516 54216 37657 54244
rect 37516 54204 37522 54216
rect 37645 54213 37657 54216
rect 37691 54213 37703 54247
rect 38378 54244 38384 54256
rect 38339 54216 38384 54244
rect 37645 54207 37703 54213
rect 38378 54204 38384 54216
rect 38436 54204 38442 54256
rect 38562 54244 38568 54256
rect 38523 54216 38568 54244
rect 38562 54204 38568 54216
rect 38620 54204 38626 54256
rect 39761 54247 39819 54253
rect 39761 54213 39773 54247
rect 39807 54244 39819 54247
rect 39942 54244 39948 54256
rect 39807 54216 39948 54244
rect 39807 54213 39819 54216
rect 39761 54207 39819 54213
rect 39942 54204 39948 54216
rect 40000 54204 40006 54256
rect 42076 54191 42104 54272
rect 32217 54179 32275 54185
rect 32217 54145 32229 54179
rect 32263 54145 32275 54179
rect 32217 54139 32275 54145
rect 32398 54136 32404 54188
rect 32456 54176 32462 54188
rect 32493 54179 32551 54185
rect 32493 54176 32505 54179
rect 32456 54148 32505 54176
rect 32456 54136 32462 54148
rect 32493 54145 32505 54148
rect 32539 54145 32551 54179
rect 32493 54139 32551 54145
rect 33873 54179 33931 54185
rect 33873 54145 33885 54179
rect 33919 54176 33931 54179
rect 34238 54176 34244 54188
rect 33919 54148 34244 54176
rect 33919 54145 33931 54148
rect 33873 54139 33931 54145
rect 34238 54136 34244 54148
rect 34296 54136 34302 54188
rect 34698 54176 34704 54188
rect 34659 54148 34704 54176
rect 34698 54136 34704 54148
rect 34756 54136 34762 54188
rect 34974 54176 34980 54188
rect 34935 54148 34980 54176
rect 34974 54136 34980 54148
rect 35032 54136 35038 54188
rect 35618 54176 35624 54188
rect 35579 54148 35624 54176
rect 35618 54136 35624 54148
rect 35676 54136 35682 54188
rect 36078 54176 36084 54188
rect 36039 54148 36084 54176
rect 36078 54136 36084 54148
rect 36136 54136 36142 54188
rect 36354 54136 36360 54188
rect 36412 54176 36418 54188
rect 37001 54179 37059 54185
rect 37001 54176 37013 54179
rect 36412 54148 37013 54176
rect 36412 54136 36418 54148
rect 37001 54145 37013 54148
rect 37047 54145 37059 54179
rect 37001 54139 37059 54145
rect 39485 54179 39543 54185
rect 39485 54145 39497 54179
rect 39531 54176 39543 54179
rect 39666 54176 39672 54188
rect 39531 54148 39672 54176
rect 39531 54145 39543 54148
rect 39485 54139 39543 54145
rect 39666 54136 39672 54148
rect 39724 54136 39730 54188
rect 40310 54136 40316 54188
rect 40368 54176 40374 54188
rect 40770 54176 40776 54188
rect 40368 54148 40776 54176
rect 40368 54136 40374 54148
rect 40770 54136 40776 54148
rect 40828 54176 40834 54188
rect 40957 54179 41015 54185
rect 40957 54176 40969 54179
rect 40828 54148 40969 54176
rect 40828 54136 40834 54148
rect 40957 54145 40969 54148
rect 41003 54145 41015 54179
rect 40957 54139 41015 54145
rect 41690 54136 41696 54188
rect 41748 54176 41754 54188
rect 42071 54185 42129 54191
rect 41973 54179 42031 54185
rect 41973 54176 41985 54179
rect 41748 54148 41985 54176
rect 41748 54136 41754 54148
rect 41973 54145 41985 54148
rect 42019 54145 42031 54179
rect 42071 54151 42083 54185
rect 42117 54151 42129 54185
rect 42071 54145 42129 54151
rect 42189 54179 42247 54185
rect 42189 54145 42201 54179
rect 42235 54176 42247 54179
rect 42426 54176 42432 54188
rect 42235 54148 42432 54176
rect 42235 54145 42247 54148
rect 41973 54139 42031 54145
rect 42189 54139 42247 54145
rect 42426 54136 42432 54148
rect 42484 54136 42490 54188
rect 30944 54108 30972 54136
rect 32033 54111 32091 54117
rect 32033 54108 32045 54111
rect 29656 54080 32045 54108
rect 32033 54077 32045 54080
rect 32079 54077 32091 54111
rect 32033 54071 32091 54077
rect 33965 54111 34023 54117
rect 33965 54077 33977 54111
rect 34011 54108 34023 54111
rect 34517 54111 34575 54117
rect 34517 54108 34529 54111
rect 34011 54080 34529 54108
rect 34011 54077 34023 54080
rect 33965 54071 34023 54077
rect 34517 54077 34529 54080
rect 34563 54077 34575 54111
rect 34882 54108 34888 54120
rect 34843 54080 34888 54108
rect 34517 54071 34575 54077
rect 34882 54068 34888 54080
rect 34940 54068 34946 54120
rect 40218 54108 40224 54120
rect 39776 54080 40224 54108
rect 26418 54000 26424 54052
rect 26476 54040 26482 54052
rect 27338 54040 27344 54052
rect 26476 54012 27344 54040
rect 26476 54000 26482 54012
rect 27338 54000 27344 54012
rect 27396 54040 27402 54052
rect 28166 54040 28172 54052
rect 27396 54012 28172 54040
rect 27396 54000 27402 54012
rect 28166 54000 28172 54012
rect 28224 54000 28230 54052
rect 29362 54040 29368 54052
rect 29323 54012 29368 54040
rect 29362 54000 29368 54012
rect 29420 54000 29426 54052
rect 31205 54043 31263 54049
rect 31205 54009 31217 54043
rect 31251 54040 31263 54043
rect 31662 54040 31668 54052
rect 31251 54012 31668 54040
rect 31251 54009 31263 54012
rect 31205 54003 31263 54009
rect 31662 54000 31668 54012
rect 31720 54000 31726 54052
rect 39776 54049 39804 54080
rect 40218 54068 40224 54080
rect 40276 54068 40282 54120
rect 39761 54043 39819 54049
rect 39761 54009 39773 54043
rect 39807 54009 39819 54043
rect 39761 54003 39819 54009
rect 28537 53975 28595 53981
rect 28537 53941 28549 53975
rect 28583 53972 28595 53975
rect 32030 53972 32036 53984
rect 28583 53944 32036 53972
rect 28583 53941 28595 53944
rect 28537 53935 28595 53941
rect 32030 53932 32036 53944
rect 32088 53932 32094 53984
rect 40034 53932 40040 53984
rect 40092 53972 40098 53984
rect 40221 53975 40279 53981
rect 40221 53972 40233 53975
rect 40092 53944 40233 53972
rect 40092 53932 40098 53944
rect 40221 53941 40233 53944
rect 40267 53941 40279 53975
rect 40221 53935 40279 53941
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 28166 53768 28172 53780
rect 28127 53740 28172 53768
rect 28166 53728 28172 53740
rect 28224 53728 28230 53780
rect 29178 53728 29184 53780
rect 29236 53768 29242 53780
rect 29273 53771 29331 53777
rect 29273 53768 29285 53771
rect 29236 53740 29285 53768
rect 29236 53728 29242 53740
rect 29273 53737 29285 53740
rect 29319 53737 29331 53771
rect 29273 53731 29331 53737
rect 29914 53728 29920 53780
rect 29972 53768 29978 53780
rect 30009 53771 30067 53777
rect 30009 53768 30021 53771
rect 29972 53740 30021 53768
rect 29972 53728 29978 53740
rect 30009 53737 30021 53740
rect 30055 53737 30067 53771
rect 30009 53731 30067 53737
rect 32677 53771 32735 53777
rect 32677 53737 32689 53771
rect 32723 53768 32735 53771
rect 32766 53768 32772 53780
rect 32723 53740 32772 53768
rect 32723 53737 32735 53740
rect 32677 53731 32735 53737
rect 32766 53728 32772 53740
rect 32824 53728 32830 53780
rect 33594 53768 33600 53780
rect 33555 53740 33600 53768
rect 33594 53728 33600 53740
rect 33652 53728 33658 53780
rect 33781 53771 33839 53777
rect 33781 53737 33793 53771
rect 33827 53768 33839 53771
rect 34422 53768 34428 53780
rect 33827 53740 34428 53768
rect 33827 53737 33839 53740
rect 33781 53731 33839 53737
rect 28813 53635 28871 53641
rect 28813 53601 28825 53635
rect 28859 53632 28871 53635
rect 33796 53632 33824 53731
rect 34422 53728 34428 53740
rect 34480 53728 34486 53780
rect 35618 53728 35624 53780
rect 35676 53768 35682 53780
rect 35713 53771 35771 53777
rect 35713 53768 35725 53771
rect 35676 53740 35725 53768
rect 35676 53728 35682 53740
rect 35713 53737 35725 53740
rect 35759 53737 35771 53771
rect 35713 53731 35771 53737
rect 35894 53728 35900 53780
rect 35952 53768 35958 53780
rect 36817 53771 36875 53777
rect 36817 53768 36829 53771
rect 35952 53740 36829 53768
rect 35952 53728 35958 53740
rect 36817 53737 36829 53740
rect 36863 53737 36875 53771
rect 36817 53731 36875 53737
rect 37734 53728 37740 53780
rect 37792 53768 37798 53780
rect 37829 53771 37887 53777
rect 37829 53768 37841 53771
rect 37792 53740 37841 53768
rect 37792 53728 37798 53740
rect 37829 53737 37841 53740
rect 37875 53737 37887 53771
rect 37829 53731 37887 53737
rect 38838 53728 38844 53780
rect 38896 53768 38902 53780
rect 38933 53771 38991 53777
rect 38933 53768 38945 53771
rect 38896 53740 38945 53768
rect 38896 53728 38902 53740
rect 38933 53737 38945 53740
rect 38979 53737 38991 53771
rect 38933 53731 38991 53737
rect 39669 53771 39727 53777
rect 39669 53737 39681 53771
rect 39715 53768 39727 53771
rect 39850 53768 39856 53780
rect 39715 53740 39856 53768
rect 39715 53737 39727 53740
rect 39669 53731 39727 53737
rect 39850 53728 39856 53740
rect 39908 53728 39914 53780
rect 39942 53728 39948 53780
rect 40000 53768 40006 53780
rect 40221 53771 40279 53777
rect 40221 53768 40233 53771
rect 40000 53740 40233 53768
rect 40000 53728 40006 53740
rect 40221 53737 40233 53740
rect 40267 53737 40279 53771
rect 40770 53768 40776 53780
rect 40731 53740 40776 53768
rect 40221 53731 40279 53737
rect 36357 53703 36415 53709
rect 36357 53669 36369 53703
rect 36403 53700 36415 53703
rect 37458 53700 37464 53712
rect 36403 53672 37464 53700
rect 36403 53669 36415 53672
rect 36357 53663 36415 53669
rect 37458 53660 37464 53672
rect 37516 53660 37522 53712
rect 40236 53700 40264 53731
rect 40770 53728 40776 53740
rect 40828 53728 40834 53780
rect 41417 53771 41475 53777
rect 41417 53768 41429 53771
rect 41340 53740 41429 53768
rect 41340 53700 41368 53740
rect 41417 53737 41429 53740
rect 41463 53768 41475 53771
rect 42702 53768 42708 53780
rect 41463 53740 42708 53768
rect 41463 53737 41475 53740
rect 41417 53731 41475 53737
rect 42702 53728 42708 53740
rect 42760 53728 42766 53780
rect 40236 53672 41368 53700
rect 28859 53604 29408 53632
rect 28859 53601 28871 53604
rect 28813 53595 28871 53601
rect 29380 53576 29408 53604
rect 33060 53604 33824 53632
rect 29270 53564 29276 53576
rect 29231 53536 29276 53564
rect 29270 53524 29276 53536
rect 29328 53524 29334 53576
rect 29362 53524 29368 53576
rect 29420 53564 29426 53576
rect 29457 53567 29515 53573
rect 29457 53564 29469 53567
rect 29420 53536 29469 53564
rect 29420 53524 29426 53536
rect 29457 53533 29469 53536
rect 29503 53564 29515 53567
rect 30282 53564 30288 53576
rect 29503 53536 30288 53564
rect 29503 53533 29515 53536
rect 29457 53527 29515 53533
rect 30282 53524 30288 53536
rect 30340 53524 30346 53576
rect 31386 53524 31392 53576
rect 31444 53564 31450 53576
rect 33060 53573 33088 53604
rect 32861 53567 32919 53573
rect 32861 53564 32873 53567
rect 31444 53536 32873 53564
rect 31444 53524 31450 53536
rect 32861 53533 32873 53536
rect 32907 53533 32919 53567
rect 32861 53527 32919 53533
rect 33045 53567 33103 53573
rect 33045 53533 33057 53567
rect 33091 53533 33103 53567
rect 33045 53527 33103 53533
rect 31389 53431 31447 53437
rect 31389 53397 31401 53431
rect 31435 53428 31447 53431
rect 31938 53428 31944 53440
rect 31435 53400 31944 53428
rect 31435 53397 31447 53400
rect 31389 53391 31447 53397
rect 31938 53388 31944 53400
rect 31996 53388 32002 53440
rect 32876 53428 32904 53527
rect 33134 53524 33140 53576
rect 33192 53564 33198 53576
rect 35161 53567 35219 53573
rect 33192 53536 33237 53564
rect 33192 53524 33198 53536
rect 35161 53533 35173 53567
rect 35207 53564 35219 53567
rect 36078 53564 36084 53576
rect 35207 53536 36084 53564
rect 35207 53533 35219 53536
rect 35161 53527 35219 53533
rect 36078 53524 36084 53536
rect 36136 53524 36142 53576
rect 39761 53567 39819 53573
rect 39761 53533 39773 53567
rect 39807 53564 39819 53567
rect 39942 53564 39948 53576
rect 39807 53536 39948 53564
rect 39807 53533 39819 53536
rect 39761 53527 39819 53533
rect 39942 53524 39948 53536
rect 40000 53524 40006 53576
rect 33152 53496 33180 53524
rect 33760 53499 33818 53505
rect 33760 53496 33772 53499
rect 33152 53468 33772 53496
rect 33760 53465 33772 53468
rect 33806 53465 33818 53499
rect 33760 53459 33818 53465
rect 33965 53499 34023 53505
rect 33965 53465 33977 53499
rect 34011 53496 34023 53499
rect 34146 53496 34152 53508
rect 34011 53468 34152 53496
rect 34011 53465 34023 53468
rect 33965 53459 34023 53465
rect 33980 53428 34008 53459
rect 34146 53456 34152 53468
rect 34204 53456 34210 53508
rect 32876 53400 34008 53428
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 30282 53224 30288 53236
rect 30195 53196 30288 53224
rect 30282 53184 30288 53196
rect 30340 53224 30346 53236
rect 31938 53224 31944 53236
rect 30340 53196 31944 53224
rect 30340 53184 30346 53196
rect 31938 53184 31944 53196
rect 31996 53224 32002 53236
rect 33689 53227 33747 53233
rect 33689 53224 33701 53227
rect 31996 53196 33701 53224
rect 31996 53184 32002 53196
rect 33689 53193 33701 53196
rect 33735 53224 33747 53227
rect 35618 53224 35624 53236
rect 33735 53196 35624 53224
rect 33735 53193 33747 53196
rect 33689 53187 33747 53193
rect 35618 53184 35624 53196
rect 35676 53184 35682 53236
rect 38654 53184 38660 53236
rect 38712 53224 38718 53236
rect 39025 53227 39083 53233
rect 39025 53224 39037 53227
rect 38712 53196 39037 53224
rect 38712 53184 38718 53196
rect 39025 53193 39037 53196
rect 39071 53193 39083 53227
rect 39942 53224 39948 53236
rect 39903 53196 39948 53224
rect 39025 53187 39083 53193
rect 39942 53184 39948 53196
rect 40000 53224 40006 53236
rect 40957 53227 41015 53233
rect 40957 53224 40969 53227
rect 40000 53196 40969 53224
rect 40000 53184 40006 53196
rect 40957 53193 40969 53196
rect 41003 53193 41015 53227
rect 40957 53187 41015 53193
rect 33137 53159 33195 53165
rect 33137 53125 33149 53159
rect 33183 53156 33195 53159
rect 33778 53156 33784 53168
rect 33183 53128 33784 53156
rect 33183 53125 33195 53128
rect 33137 53119 33195 53125
rect 33778 53116 33784 53128
rect 33836 53116 33842 53168
rect 35897 53159 35955 53165
rect 35897 53125 35909 53159
rect 35943 53156 35955 53159
rect 36446 53156 36452 53168
rect 35943 53128 36452 53156
rect 35943 53125 35955 53128
rect 35897 53119 35955 53125
rect 36446 53116 36452 53128
rect 36504 53116 36510 53168
rect 38565 53159 38623 53165
rect 38565 53125 38577 53159
rect 38611 53156 38623 53159
rect 39960 53156 39988 53184
rect 38611 53128 39988 53156
rect 38611 53125 38623 53128
rect 38565 53119 38623 53125
rect 29454 53048 29460 53100
rect 29512 53088 29518 53100
rect 29549 53091 29607 53097
rect 29549 53088 29561 53091
rect 29512 53060 29561 53088
rect 29512 53048 29518 53060
rect 29549 53057 29561 53060
rect 29595 53057 29607 53091
rect 29549 53051 29607 53057
rect 36078 53048 36084 53100
rect 36136 53088 36142 53100
rect 36136 53060 36181 53088
rect 36136 53048 36142 53060
rect 34514 53020 34520 53032
rect 34475 52992 34520 53020
rect 34514 52980 34520 52992
rect 34572 52980 34578 53032
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 29362 52680 29368 52692
rect 29323 52652 29368 52680
rect 29362 52640 29368 52652
rect 29420 52640 29426 52692
rect 35069 52683 35127 52689
rect 35069 52649 35081 52683
rect 35115 52680 35127 52683
rect 35618 52680 35624 52692
rect 35115 52652 35624 52680
rect 35115 52649 35127 52652
rect 35069 52643 35127 52649
rect 35618 52640 35624 52652
rect 35676 52640 35682 52692
rect 36081 52683 36139 52689
rect 36081 52649 36093 52683
rect 36127 52680 36139 52683
rect 36170 52680 36176 52692
rect 36127 52652 36176 52680
rect 36127 52649 36139 52652
rect 36081 52643 36139 52649
rect 36170 52640 36176 52652
rect 36228 52640 36234 52692
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 26418 8072 26424 8084
rect 26379 8044 26424 8072
rect 26418 8032 26424 8044
rect 26476 8032 26482 8084
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 24946 7420 24952 7472
rect 25004 7460 25010 7472
rect 25961 7463 26019 7469
rect 25961 7460 25973 7463
rect 25004 7432 25973 7460
rect 25004 7420 25010 7432
rect 25961 7429 25973 7432
rect 26007 7429 26019 7463
rect 25961 7423 26019 7429
rect 29641 7395 29699 7401
rect 29641 7361 29653 7395
rect 29687 7392 29699 7395
rect 30282 7392 30288 7404
rect 29687 7364 30288 7392
rect 29687 7361 29699 7364
rect 29641 7355 29699 7361
rect 30282 7352 30288 7364
rect 30340 7352 30346 7404
rect 22554 7284 22560 7336
rect 22612 7324 22618 7336
rect 25777 7327 25835 7333
rect 25777 7324 25789 7327
rect 22612 7296 25789 7324
rect 22612 7284 22618 7296
rect 25777 7293 25789 7296
rect 25823 7293 25835 7327
rect 26786 7324 26792 7336
rect 26747 7296 26792 7324
rect 25777 7287 25835 7293
rect 26786 7284 26792 7296
rect 26844 7284 26850 7336
rect 26694 7148 26700 7200
rect 26752 7188 26758 7200
rect 28077 7191 28135 7197
rect 28077 7188 28089 7191
rect 26752 7160 28089 7188
rect 26752 7148 26758 7160
rect 28077 7157 28089 7160
rect 28123 7157 28135 7191
rect 29730 7188 29736 7200
rect 29691 7160 29736 7188
rect 28077 7151 28135 7157
rect 29730 7148 29736 7160
rect 29788 7148 29794 7200
rect 30374 7188 30380 7200
rect 30335 7160 30380 7188
rect 30374 7148 30380 7160
rect 30432 7148 30438 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 25590 6808 25596 6860
rect 25648 6848 25654 6860
rect 27985 6851 28043 6857
rect 27985 6848 27997 6851
rect 25648 6820 27997 6848
rect 25648 6808 25654 6820
rect 27985 6817 27997 6820
rect 28031 6817 28043 6851
rect 28626 6848 28632 6860
rect 28587 6820 28632 6848
rect 27985 6811 28043 6817
rect 28626 6808 28632 6820
rect 28684 6808 28690 6860
rect 25961 6783 26019 6789
rect 25961 6749 25973 6783
rect 26007 6780 26019 6783
rect 26007 6752 26234 6780
rect 26007 6749 26019 6752
rect 25961 6743 26019 6749
rect 26206 6712 26234 6752
rect 26602 6740 26608 6792
rect 26660 6780 26666 6792
rect 27341 6783 27399 6789
rect 27341 6780 27353 6783
rect 26660 6752 27353 6780
rect 26660 6740 26666 6752
rect 27341 6749 27353 6752
rect 27387 6749 27399 6783
rect 27341 6743 27399 6749
rect 29546 6740 29552 6792
rect 29604 6780 29610 6792
rect 30285 6783 30343 6789
rect 30285 6780 30297 6783
rect 29604 6752 30297 6780
rect 29604 6740 29610 6752
rect 30285 6749 30297 6752
rect 30331 6749 30343 6783
rect 31018 6780 31024 6792
rect 30979 6752 31024 6780
rect 30285 6743 30343 6749
rect 31018 6740 31024 6752
rect 31076 6740 31082 6792
rect 31754 6740 31760 6792
rect 31812 6780 31818 6792
rect 32125 6783 32183 6789
rect 32125 6780 32137 6783
rect 31812 6752 32137 6780
rect 31812 6740 31818 6752
rect 32125 6749 32137 6752
rect 32171 6749 32183 6783
rect 32125 6743 32183 6749
rect 26510 6712 26516 6724
rect 26206 6684 26516 6712
rect 26510 6672 26516 6684
rect 26568 6712 26574 6724
rect 28166 6712 28172 6724
rect 26568 6684 28028 6712
rect 28127 6684 28172 6712
rect 26568 6672 26574 6684
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 25869 6647 25927 6653
rect 25869 6644 25881 6647
rect 24912 6616 25881 6644
rect 24912 6604 24918 6616
rect 25869 6613 25881 6616
rect 25915 6613 25927 6647
rect 25869 6607 25927 6613
rect 26878 6604 26884 6656
rect 26936 6644 26942 6656
rect 27433 6647 27491 6653
rect 27433 6644 27445 6647
rect 26936 6616 27445 6644
rect 26936 6604 26942 6616
rect 27433 6613 27445 6616
rect 27479 6613 27491 6647
rect 28000 6644 28028 6684
rect 28166 6672 28172 6684
rect 28224 6672 28230 6724
rect 30374 6644 30380 6656
rect 28000 6616 30380 6644
rect 27433 6607 27491 6613
rect 30374 6604 30380 6616
rect 30432 6604 30438 6656
rect 32214 6644 32220 6656
rect 32175 6616 32220 6644
rect 32214 6604 32220 6616
rect 32272 6604 32278 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 26145 6375 26203 6381
rect 26145 6341 26157 6375
rect 26191 6372 26203 6375
rect 26881 6375 26939 6381
rect 26881 6372 26893 6375
rect 26191 6344 26893 6372
rect 26191 6341 26203 6344
rect 26145 6335 26203 6341
rect 26881 6341 26893 6344
rect 26927 6341 26939 6375
rect 29730 6372 29736 6384
rect 29691 6344 29736 6372
rect 26881 6335 26939 6341
rect 29730 6332 29736 6344
rect 29788 6332 29794 6384
rect 35621 6375 35679 6381
rect 35621 6341 35633 6375
rect 35667 6372 35679 6375
rect 38194 6372 38200 6384
rect 35667 6344 38200 6372
rect 35667 6341 35679 6344
rect 35621 6335 35679 6341
rect 38194 6332 38200 6344
rect 38252 6332 38258 6384
rect 24486 6264 24492 6316
rect 24544 6304 24550 6316
rect 26053 6307 26111 6313
rect 26053 6304 26065 6307
rect 24544 6276 26065 6304
rect 24544 6264 24550 6276
rect 26053 6273 26065 6276
rect 26099 6304 26111 6307
rect 26602 6304 26608 6316
rect 26099 6276 26608 6304
rect 26099 6273 26111 6276
rect 26053 6267 26111 6273
rect 26602 6264 26608 6276
rect 26660 6264 26666 6316
rect 29546 6304 29552 6316
rect 29507 6276 29552 6304
rect 29546 6264 29552 6276
rect 29604 6264 29610 6316
rect 31849 6307 31907 6313
rect 31849 6273 31861 6307
rect 31895 6273 31907 6307
rect 31849 6267 31907 6273
rect 26234 6196 26240 6248
rect 26292 6236 26298 6248
rect 26697 6239 26755 6245
rect 26697 6236 26709 6239
rect 26292 6208 26709 6236
rect 26292 6196 26298 6208
rect 26697 6205 26709 6208
rect 26743 6205 26755 6239
rect 27890 6236 27896 6248
rect 27851 6208 27896 6236
rect 26697 6199 26755 6205
rect 27890 6196 27896 6208
rect 27948 6196 27954 6248
rect 30190 6236 30196 6248
rect 30151 6208 30196 6236
rect 30190 6196 30196 6208
rect 30248 6196 30254 6248
rect 30282 6196 30288 6248
rect 30340 6236 30346 6248
rect 31864 6236 31892 6267
rect 34422 6236 34428 6248
rect 30340 6208 31892 6236
rect 34383 6208 34428 6236
rect 30340 6196 30346 6208
rect 34422 6196 34428 6208
rect 34480 6196 34486 6248
rect 35805 6239 35863 6245
rect 35805 6205 35817 6239
rect 35851 6236 35863 6239
rect 37918 6236 37924 6248
rect 35851 6208 37924 6236
rect 35851 6205 35863 6208
rect 35805 6199 35863 6205
rect 37918 6196 37924 6208
rect 37976 6196 37982 6248
rect 23934 6060 23940 6112
rect 23992 6100 23998 6112
rect 24029 6103 24087 6109
rect 24029 6100 24041 6103
rect 23992 6072 24041 6100
rect 23992 6060 23998 6072
rect 24029 6069 24041 6072
rect 24075 6069 24087 6103
rect 24029 6063 24087 6069
rect 24670 6060 24676 6112
rect 24728 6100 24734 6112
rect 25409 6103 25467 6109
rect 25409 6100 25421 6103
rect 24728 6072 25421 6100
rect 24728 6060 24734 6072
rect 25409 6069 25421 6072
rect 25455 6069 25467 6103
rect 25409 6063 25467 6069
rect 31202 6060 31208 6112
rect 31260 6100 31266 6112
rect 31941 6103 31999 6109
rect 31941 6100 31953 6103
rect 31260 6072 31953 6100
rect 31260 6060 31266 6072
rect 31941 6069 31953 6072
rect 31987 6069 31999 6103
rect 33042 6100 33048 6112
rect 33003 6072 33048 6100
rect 31941 6063 31999 6069
rect 33042 6060 33048 6072
rect 33100 6060 33106 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 24670 5760 24676 5772
rect 24631 5732 24676 5760
rect 24670 5720 24676 5732
rect 24728 5720 24734 5772
rect 24854 5760 24860 5772
rect 24815 5732 24860 5760
rect 24854 5720 24860 5732
rect 24912 5720 24918 5772
rect 26142 5760 26148 5772
rect 26103 5732 26148 5760
rect 26142 5720 26148 5732
rect 26200 5720 26206 5772
rect 28074 5760 28080 5772
rect 28035 5732 28080 5760
rect 28074 5720 28080 5732
rect 28132 5720 28138 5772
rect 30098 5720 30104 5772
rect 30156 5760 30162 5772
rect 30282 5760 30288 5772
rect 30156 5732 30288 5760
rect 30156 5720 30162 5732
rect 30282 5720 30288 5732
rect 30340 5720 30346 5772
rect 31018 5760 31024 5772
rect 30979 5732 31024 5760
rect 31018 5720 31024 5732
rect 31076 5720 31082 5772
rect 31202 5760 31208 5772
rect 31163 5732 31208 5760
rect 31202 5720 31208 5732
rect 31260 5720 31266 5772
rect 31662 5760 31668 5772
rect 31623 5732 31668 5760
rect 31662 5720 31668 5732
rect 31720 5720 31726 5772
rect 23106 5652 23112 5704
rect 23164 5692 23170 5704
rect 23201 5695 23259 5701
rect 23201 5692 23213 5695
rect 23164 5664 23213 5692
rect 23164 5652 23170 5664
rect 23201 5661 23213 5664
rect 23247 5661 23259 5695
rect 23201 5655 23259 5661
rect 24213 5695 24271 5701
rect 24213 5661 24225 5695
rect 24259 5692 24271 5695
rect 24486 5692 24492 5704
rect 24259 5664 24492 5692
rect 24259 5661 24271 5664
rect 24213 5655 24271 5661
rect 24486 5652 24492 5664
rect 24544 5652 24550 5704
rect 26050 5652 26056 5704
rect 26108 5692 26114 5704
rect 26510 5692 26516 5704
rect 26108 5664 26516 5692
rect 26108 5652 26114 5664
rect 26510 5652 26516 5664
rect 26568 5652 26574 5704
rect 27522 5692 27528 5704
rect 27483 5664 27528 5692
rect 27522 5652 27528 5664
rect 27580 5652 27586 5704
rect 30009 5695 30067 5701
rect 30009 5661 30021 5695
rect 30055 5692 30067 5695
rect 30374 5692 30380 5704
rect 30055 5664 30380 5692
rect 30055 5661 30067 5664
rect 30009 5655 30067 5661
rect 30374 5652 30380 5664
rect 30432 5692 30438 5704
rect 30432 5664 31064 5692
rect 30432 5652 30438 5664
rect 31036 5636 31064 5664
rect 33134 5652 33140 5704
rect 33192 5692 33198 5704
rect 33321 5695 33379 5701
rect 33321 5692 33333 5695
rect 33192 5664 33333 5692
rect 33192 5652 33198 5664
rect 33321 5661 33333 5664
rect 33367 5661 33379 5695
rect 33321 5655 33379 5661
rect 34149 5695 34207 5701
rect 34149 5661 34161 5695
rect 34195 5692 34207 5695
rect 35161 5695 35219 5701
rect 35161 5692 35173 5695
rect 34195 5664 35173 5692
rect 34195 5661 34207 5664
rect 34149 5655 34207 5661
rect 35161 5661 35173 5664
rect 35207 5692 35219 5695
rect 35342 5692 35348 5704
rect 35207 5664 35348 5692
rect 35207 5661 35219 5664
rect 35161 5655 35219 5661
rect 26970 5584 26976 5636
rect 27028 5624 27034 5636
rect 27709 5627 27767 5633
rect 27709 5624 27721 5627
rect 27028 5596 27721 5624
rect 27028 5584 27034 5596
rect 27709 5593 27721 5596
rect 27755 5593 27767 5627
rect 27709 5587 27767 5593
rect 31018 5584 31024 5636
rect 31076 5584 31082 5636
rect 31754 5584 31760 5636
rect 31812 5624 31818 5636
rect 34164 5624 34192 5655
rect 35342 5652 35348 5664
rect 35400 5652 35406 5704
rect 31812 5596 34192 5624
rect 31812 5584 31818 5596
rect 24118 5556 24124 5568
rect 24079 5528 24124 5556
rect 24118 5516 24124 5528
rect 24176 5516 24182 5568
rect 33226 5516 33232 5568
rect 33284 5556 33290 5568
rect 34057 5559 34115 5565
rect 34057 5556 34069 5559
rect 33284 5528 34069 5556
rect 33284 5516 33290 5528
rect 34057 5525 34069 5528
rect 34103 5525 34115 5559
rect 34057 5519 34115 5525
rect 34790 5516 34796 5568
rect 34848 5556 34854 5568
rect 35069 5559 35127 5565
rect 35069 5556 35081 5559
rect 34848 5528 35081 5556
rect 34848 5516 34854 5528
rect 35069 5525 35081 5528
rect 35115 5525 35127 5559
rect 35069 5519 35127 5525
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 25225 5355 25283 5361
rect 25225 5321 25237 5355
rect 25271 5352 25283 5355
rect 26970 5352 26976 5364
rect 25271 5324 26976 5352
rect 25271 5321 25283 5324
rect 25225 5315 25283 5321
rect 26970 5312 26976 5324
rect 27028 5312 27034 5364
rect 22925 5287 22983 5293
rect 22925 5253 22937 5287
rect 22971 5284 22983 5287
rect 24118 5284 24124 5296
rect 22971 5256 24124 5284
rect 22971 5253 22983 5256
rect 22925 5247 22983 5253
rect 24118 5244 24124 5256
rect 24176 5244 24182 5296
rect 26878 5284 26884 5296
rect 26839 5256 26884 5284
rect 26878 5244 26884 5256
rect 26936 5244 26942 5296
rect 34790 5284 34796 5296
rect 34751 5256 34796 5284
rect 34790 5244 34796 5256
rect 34848 5244 34854 5296
rect 24486 5176 24492 5228
rect 24544 5216 24550 5228
rect 25133 5219 25191 5225
rect 25133 5216 25145 5219
rect 24544 5188 25145 5216
rect 24544 5176 24550 5188
rect 25133 5185 25145 5188
rect 25179 5216 25191 5219
rect 25777 5219 25835 5225
rect 25179 5188 25544 5216
rect 25179 5185 25191 5188
rect 25133 5179 25191 5185
rect 22278 5108 22284 5160
rect 22336 5148 22342 5160
rect 22741 5151 22799 5157
rect 22741 5148 22753 5151
rect 22336 5120 22753 5148
rect 22336 5108 22342 5120
rect 22741 5117 22753 5120
rect 22787 5117 22799 5151
rect 22741 5111 22799 5117
rect 24581 5151 24639 5157
rect 24581 5117 24593 5151
rect 24627 5148 24639 5151
rect 25406 5148 25412 5160
rect 24627 5120 25412 5148
rect 24627 5117 24639 5120
rect 24581 5111 24639 5117
rect 25406 5108 25412 5120
rect 25464 5108 25470 5160
rect 25516 5148 25544 5188
rect 25777 5185 25789 5219
rect 25823 5216 25835 5219
rect 26050 5216 26056 5228
rect 25823 5188 26056 5216
rect 25823 5185 25835 5188
rect 25777 5179 25835 5185
rect 26050 5176 26056 5188
rect 26108 5176 26114 5228
rect 26694 5216 26700 5228
rect 26655 5188 26700 5216
rect 26694 5176 26700 5188
rect 26752 5176 26758 5228
rect 25961 5151 26019 5157
rect 25961 5148 25973 5151
rect 25516 5120 25973 5148
rect 25961 5117 25973 5120
rect 26007 5117 26019 5151
rect 28350 5148 28356 5160
rect 28311 5120 28356 5148
rect 25961 5111 26019 5117
rect 28350 5108 28356 5120
rect 28408 5108 28414 5160
rect 29641 5151 29699 5157
rect 29641 5117 29653 5151
rect 29687 5148 29699 5151
rect 30101 5151 30159 5157
rect 30101 5148 30113 5151
rect 29687 5120 30113 5148
rect 29687 5117 29699 5120
rect 29641 5111 29699 5117
rect 30101 5117 30113 5120
rect 30147 5117 30159 5151
rect 30282 5148 30288 5160
rect 30243 5120 30288 5148
rect 30101 5111 30159 5117
rect 30282 5108 30288 5120
rect 30340 5108 30346 5160
rect 30558 5148 30564 5160
rect 30519 5120 30564 5148
rect 30558 5108 30564 5120
rect 30616 5108 30622 5160
rect 33318 5148 33324 5160
rect 33279 5120 33324 5148
rect 33318 5108 33324 5120
rect 33376 5108 33382 5160
rect 34977 5151 35035 5157
rect 34977 5117 34989 5151
rect 35023 5148 35035 5151
rect 35437 5151 35495 5157
rect 35437 5148 35449 5151
rect 35023 5120 35449 5148
rect 35023 5117 35035 5120
rect 34977 5111 35035 5117
rect 35437 5117 35449 5120
rect 35483 5117 35495 5151
rect 35437 5111 35495 5117
rect 22281 5015 22339 5021
rect 22281 4981 22293 5015
rect 22327 5012 22339 5015
rect 22830 5012 22836 5024
rect 22327 4984 22836 5012
rect 22327 4981 22339 4984
rect 22281 4975 22339 4981
rect 22830 4972 22836 4984
rect 22888 4972 22894 5024
rect 31018 4972 31024 5024
rect 31076 5012 31082 5024
rect 32401 5015 32459 5021
rect 32401 5012 32413 5015
rect 31076 4984 32413 5012
rect 31076 4972 31082 4984
rect 32401 4981 32413 4984
rect 32447 4981 32459 5015
rect 32401 4975 32459 4981
rect 35894 4972 35900 5024
rect 35952 5012 35958 5024
rect 36081 5015 36139 5021
rect 36081 5012 36093 5015
rect 35952 4984 36093 5012
rect 35952 4972 35958 4984
rect 36081 4981 36093 4984
rect 36127 4981 36139 5015
rect 36081 4975 36139 4981
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 22554 4808 22560 4820
rect 22515 4780 22560 4808
rect 22554 4768 22560 4780
rect 22612 4768 22618 4820
rect 27522 4808 27528 4820
rect 27483 4780 27528 4808
rect 27522 4768 27528 4780
rect 27580 4768 27586 4820
rect 21913 4743 21971 4749
rect 21913 4709 21925 4743
rect 21959 4740 21971 4743
rect 23382 4740 23388 4752
rect 21959 4712 23388 4740
rect 21959 4709 21971 4712
rect 21913 4703 21971 4709
rect 23382 4700 23388 4712
rect 23440 4700 23446 4752
rect 33134 4740 33140 4752
rect 32048 4712 33140 4740
rect 24486 4672 24492 4684
rect 23400 4644 24492 4672
rect 19334 4604 19340 4616
rect 19295 4576 19340 4604
rect 19334 4564 19340 4576
rect 19392 4564 19398 4616
rect 20346 4564 20352 4616
rect 20404 4604 20410 4616
rect 20441 4607 20499 4613
rect 20441 4604 20453 4607
rect 20404 4576 20453 4604
rect 20404 4564 20410 4576
rect 20441 4573 20453 4576
rect 20487 4573 20499 4607
rect 20441 4567 20499 4573
rect 21269 4607 21327 4613
rect 21269 4573 21281 4607
rect 21315 4604 21327 4607
rect 21726 4604 21732 4616
rect 21315 4576 21732 4604
rect 21315 4573 21327 4576
rect 21269 4567 21327 4573
rect 21726 4564 21732 4576
rect 21784 4564 21790 4616
rect 22186 4564 22192 4616
rect 22244 4604 22250 4616
rect 23400 4613 23428 4644
rect 24486 4632 24492 4644
rect 24544 4632 24550 4684
rect 30006 4672 30012 4684
rect 29967 4644 30012 4672
rect 30006 4632 30012 4644
rect 30064 4632 30070 4684
rect 31297 4675 31355 4681
rect 31297 4641 31309 4675
rect 31343 4672 31355 4675
rect 31754 4672 31760 4684
rect 31343 4644 31760 4672
rect 31343 4641 31355 4644
rect 31297 4635 31355 4641
rect 31754 4632 31760 4644
rect 31812 4632 31818 4684
rect 32048 4681 32076 4712
rect 33134 4700 33140 4712
rect 33192 4700 33198 4752
rect 37274 4700 37280 4752
rect 37332 4740 37338 4752
rect 37921 4743 37979 4749
rect 37921 4740 37933 4743
rect 37332 4712 37933 4740
rect 37332 4700 37338 4712
rect 37921 4709 37933 4712
rect 37967 4709 37979 4743
rect 37921 4703 37979 4709
rect 32033 4675 32091 4681
rect 32033 4641 32045 4675
rect 32079 4641 32091 4675
rect 32214 4672 32220 4684
rect 32175 4644 32220 4672
rect 32033 4635 32091 4641
rect 32214 4632 32220 4644
rect 32272 4632 32278 4684
rect 32766 4672 32772 4684
rect 32727 4644 32772 4672
rect 32766 4632 32772 4644
rect 32824 4632 32830 4684
rect 23385 4607 23443 4613
rect 23385 4604 23397 4607
rect 22244 4576 23397 4604
rect 22244 4564 22250 4576
rect 23385 4573 23397 4576
rect 23431 4573 23443 4607
rect 23385 4567 23443 4573
rect 24213 4607 24271 4613
rect 24213 4573 24225 4607
rect 24259 4604 24271 4607
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 24259 4576 24685 4604
rect 24259 4573 24271 4576
rect 24213 4567 24271 4573
rect 24673 4573 24685 4576
rect 24719 4573 24731 4607
rect 24673 4567 24731 4573
rect 28169 4607 28227 4613
rect 28169 4573 28181 4607
rect 28215 4604 28227 4607
rect 28629 4607 28687 4613
rect 28629 4604 28641 4607
rect 28215 4576 28641 4604
rect 28215 4573 28227 4576
rect 28169 4567 28227 4573
rect 28629 4573 28641 4576
rect 28675 4573 28687 4607
rect 31018 4604 31024 4616
rect 30979 4576 31024 4604
rect 28629 4567 28687 4573
rect 31018 4564 31024 4576
rect 31076 4564 31082 4616
rect 36814 4564 36820 4616
rect 36872 4604 36878 4616
rect 37277 4607 37335 4613
rect 36872 4576 36917 4604
rect 36872 4564 36878 4576
rect 37277 4573 37289 4607
rect 37323 4604 37335 4607
rect 37458 4604 37464 4616
rect 37323 4576 37464 4604
rect 37323 4573 37335 4576
rect 37277 4567 37335 4573
rect 37458 4564 37464 4576
rect 37516 4564 37522 4616
rect 38930 4604 38936 4616
rect 38891 4576 38936 4604
rect 38930 4564 38936 4576
rect 38988 4564 38994 4616
rect 23477 4539 23535 4545
rect 23477 4505 23489 4539
rect 23523 4536 23535 4539
rect 24857 4539 24915 4545
rect 24857 4536 24869 4539
rect 23523 4508 24869 4536
rect 23523 4505 23535 4508
rect 23477 4499 23535 4505
rect 24857 4505 24869 4508
rect 24903 4505 24915 4539
rect 24857 4499 24915 4505
rect 26513 4539 26571 4545
rect 26513 4505 26525 4539
rect 26559 4536 26571 4539
rect 27522 4536 27528 4548
rect 26559 4508 27528 4536
rect 26559 4505 26571 4508
rect 26513 4499 26571 4505
rect 27522 4496 27528 4508
rect 27580 4496 27586 4548
rect 28813 4539 28871 4545
rect 28813 4505 28825 4539
rect 28859 4536 28871 4539
rect 29454 4536 29460 4548
rect 28859 4508 29460 4536
rect 28859 4505 28871 4508
rect 28813 4499 28871 4505
rect 29454 4496 29460 4508
rect 29512 4496 29518 4548
rect 34974 4536 34980 4548
rect 34935 4508 34980 4536
rect 34974 4496 34980 4508
rect 35032 4496 35038 4548
rect 36633 4539 36691 4545
rect 36633 4505 36645 4539
rect 36679 4536 36691 4539
rect 37366 4536 37372 4548
rect 36679 4508 37372 4536
rect 36679 4505 36691 4508
rect 36633 4499 36691 4505
rect 37366 4496 37372 4508
rect 37424 4496 37430 4548
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 30101 4267 30159 4273
rect 30101 4233 30113 4267
rect 30147 4264 30159 4267
rect 30282 4264 30288 4276
rect 30147 4236 30288 4264
rect 30147 4233 30159 4236
rect 30101 4227 30159 4233
rect 30282 4224 30288 4236
rect 30340 4224 30346 4276
rect 22278 4128 22284 4140
rect 22239 4100 22284 4128
rect 22278 4088 22284 4100
rect 22336 4088 22342 4140
rect 25590 4128 25596 4140
rect 25551 4100 25596 4128
rect 25590 4088 25596 4100
rect 25648 4088 25654 4140
rect 26234 4088 26240 4140
rect 26292 4128 26298 4140
rect 29365 4131 29423 4137
rect 26292 4100 26337 4128
rect 26292 4088 26298 4100
rect 29365 4097 29377 4131
rect 29411 4128 29423 4131
rect 29546 4128 29552 4140
rect 29411 4100 29552 4128
rect 29411 4097 29423 4100
rect 29365 4091 29423 4097
rect 29546 4088 29552 4100
rect 29604 4128 29610 4140
rect 30009 4131 30067 4137
rect 30009 4128 30021 4131
rect 29604 4100 30021 4128
rect 29604 4088 29610 4100
rect 30009 4097 30021 4100
rect 30055 4128 30067 4131
rect 30098 4128 30104 4140
rect 30055 4100 30104 4128
rect 30055 4097 30067 4100
rect 30009 4091 30067 4097
rect 30098 4088 30104 4100
rect 30156 4088 30162 4140
rect 33042 4128 33048 4140
rect 33003 4100 33048 4128
rect 33042 4088 33048 4100
rect 33100 4088 33106 4140
rect 35342 4128 35348 4140
rect 35303 4100 35348 4128
rect 35342 4088 35348 4100
rect 35400 4088 35406 4140
rect 36173 4131 36231 4137
rect 36173 4097 36185 4131
rect 36219 4128 36231 4131
rect 36814 4128 36820 4140
rect 36219 4100 36820 4128
rect 36219 4097 36231 4100
rect 36173 4091 36231 4097
rect 36814 4088 36820 4100
rect 36872 4088 36878 4140
rect 19981 4063 20039 4069
rect 19981 4029 19993 4063
rect 20027 4060 20039 4063
rect 20622 4060 20628 4072
rect 20027 4032 20628 4060
rect 20027 4029 20039 4032
rect 19981 4023 20039 4029
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 22738 4060 22744 4072
rect 22699 4032 22744 4060
rect 22738 4020 22744 4032
rect 22796 4020 22802 4072
rect 22922 4060 22928 4072
rect 22883 4032 22928 4060
rect 22922 4020 22928 4032
rect 22980 4020 22986 4072
rect 24581 4063 24639 4069
rect 24581 4029 24593 4063
rect 24627 4060 24639 4063
rect 26697 4063 26755 4069
rect 24627 4032 26234 4060
rect 24627 4029 24639 4032
rect 24581 4023 24639 4029
rect 22002 3992 22008 4004
rect 20640 3964 22008 3992
rect 16298 3884 16304 3936
rect 16356 3924 16362 3936
rect 16393 3927 16451 3933
rect 16393 3924 16405 3927
rect 16356 3896 16405 3924
rect 16356 3884 16362 3896
rect 16393 3893 16405 3896
rect 16439 3893 16451 3927
rect 16393 3887 16451 3893
rect 17586 3884 17592 3936
rect 17644 3924 17650 3936
rect 17681 3927 17739 3933
rect 17681 3924 17693 3927
rect 17644 3896 17693 3924
rect 17644 3884 17650 3896
rect 17681 3893 17693 3896
rect 17727 3893 17739 3927
rect 17681 3887 17739 3893
rect 18414 3884 18420 3936
rect 18472 3924 18478 3936
rect 18509 3927 18567 3933
rect 18509 3924 18521 3927
rect 18472 3896 18521 3924
rect 18472 3884 18478 3896
rect 18509 3893 18521 3896
rect 18555 3893 18567 3927
rect 18509 3887 18567 3893
rect 19337 3927 19395 3933
rect 19337 3893 19349 3927
rect 19383 3924 19395 3927
rect 19426 3924 19432 3936
rect 19383 3896 19432 3924
rect 19383 3893 19395 3896
rect 19337 3887 19395 3893
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 20640 3933 20668 3964
rect 22002 3952 22008 3964
rect 22060 3952 22066 4004
rect 20625 3927 20683 3933
rect 20625 3893 20637 3927
rect 20671 3893 20683 3927
rect 20625 3887 20683 3893
rect 21637 3927 21695 3933
rect 21637 3893 21649 3927
rect 21683 3924 21695 3927
rect 24486 3924 24492 3936
rect 21683 3896 24492 3924
rect 21683 3893 21695 3896
rect 21637 3887 21695 3893
rect 24486 3884 24492 3896
rect 24544 3884 24550 3936
rect 26206 3924 26234 4032
rect 26697 4029 26709 4063
rect 26743 4029 26755 4063
rect 26697 4023 26755 4029
rect 26881 4063 26939 4069
rect 26881 4029 26893 4063
rect 26927 4060 26939 4063
rect 27430 4060 27436 4072
rect 26927 4032 27436 4060
rect 26927 4029 26939 4032
rect 26881 4023 26939 4029
rect 26712 3992 26740 4023
rect 27430 4020 27436 4032
rect 27488 4020 27494 4072
rect 28537 4063 28595 4069
rect 28537 4029 28549 4063
rect 28583 4060 28595 4063
rect 29730 4060 29736 4072
rect 28583 4032 29736 4060
rect 28583 4029 28595 4032
rect 28537 4023 28595 4029
rect 29730 4020 29736 4032
rect 29788 4020 29794 4072
rect 30650 4060 30656 4072
rect 30611 4032 30656 4060
rect 30650 4020 30656 4032
rect 30708 4020 30714 4072
rect 30837 4063 30895 4069
rect 30837 4029 30849 4063
rect 30883 4029 30895 4063
rect 31386 4060 31392 4072
rect 31347 4032 31392 4060
rect 30837 4023 30895 4029
rect 27982 3992 27988 4004
rect 26712 3964 27988 3992
rect 27982 3952 27988 3964
rect 28040 3952 28046 4004
rect 29457 3995 29515 4001
rect 29457 3961 29469 3995
rect 29503 3992 29515 3995
rect 30852 3992 30880 4023
rect 31386 4020 31392 4032
rect 31444 4020 31450 4072
rect 33226 4060 33232 4072
rect 33187 4032 33232 4060
rect 33226 4020 33232 4032
rect 33284 4020 33290 4072
rect 33505 4063 33563 4069
rect 33505 4029 33517 4063
rect 33551 4029 33563 4063
rect 36998 4060 37004 4072
rect 36959 4032 37004 4060
rect 33505 4023 33563 4029
rect 29503 3964 30880 3992
rect 29503 3961 29515 3964
rect 29457 3955 29515 3961
rect 33042 3952 33048 4004
rect 33100 3992 33106 4004
rect 33520 3992 33548 4023
rect 36998 4020 37004 4032
rect 37056 4020 37062 4072
rect 37182 4060 37188 4072
rect 37143 4032 37188 4060
rect 37182 4020 37188 4032
rect 37240 4020 37246 4072
rect 37461 4063 37519 4069
rect 37461 4029 37473 4063
rect 37507 4029 37519 4063
rect 37461 4023 37519 4029
rect 33100 3964 33548 3992
rect 33100 3952 33106 3964
rect 34146 3952 34152 4004
rect 34204 3992 34210 4004
rect 34204 3964 35894 3992
rect 34204 3952 34210 3964
rect 27246 3924 27252 3936
rect 26206 3896 27252 3924
rect 27246 3884 27252 3896
rect 27304 3884 27310 3936
rect 33870 3884 33876 3936
rect 33928 3924 33934 3936
rect 34974 3924 34980 3936
rect 33928 3896 34980 3924
rect 33928 3884 33934 3896
rect 34974 3884 34980 3896
rect 35032 3884 35038 3936
rect 35434 3924 35440 3936
rect 35395 3896 35440 3924
rect 35434 3884 35440 3896
rect 35492 3884 35498 3936
rect 35866 3924 35894 3964
rect 37476 3924 37504 4023
rect 39114 3952 39120 4004
rect 39172 3992 39178 4004
rect 39945 3995 40003 4001
rect 39945 3992 39957 3995
rect 39172 3964 39957 3992
rect 39172 3952 39178 3964
rect 39945 3961 39957 3964
rect 39991 3961 40003 3995
rect 39945 3955 40003 3961
rect 35866 3896 37504 3924
rect 37734 3884 37740 3936
rect 37792 3924 37798 3936
rect 39301 3927 39359 3933
rect 39301 3924 39313 3927
rect 37792 3896 39313 3924
rect 37792 3884 37798 3896
rect 39301 3893 39313 3896
rect 39347 3893 39359 3927
rect 39301 3887 39359 3893
rect 40218 3884 40224 3936
rect 40276 3924 40282 3936
rect 40957 3927 41015 3933
rect 40957 3924 40969 3927
rect 40276 3896 40969 3924
rect 40276 3884 40282 3896
rect 40957 3893 40969 3896
rect 41003 3893 41015 3927
rect 40957 3887 41015 3893
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 22738 3680 22744 3732
rect 22796 3720 22802 3732
rect 23385 3723 23443 3729
rect 23385 3720 23397 3723
rect 22796 3692 23397 3720
rect 22796 3680 22802 3692
rect 23385 3689 23397 3692
rect 23431 3689 23443 3723
rect 27430 3720 27436 3732
rect 27391 3692 27436 3720
rect 23385 3683 23443 3689
rect 27430 3680 27436 3692
rect 27488 3680 27494 3732
rect 27982 3720 27988 3732
rect 27943 3692 27988 3720
rect 27982 3680 27988 3692
rect 28040 3680 28046 3732
rect 30650 3680 30656 3732
rect 30708 3720 30714 3732
rect 31021 3723 31079 3729
rect 31021 3720 31033 3723
rect 30708 3692 31033 3720
rect 30708 3680 30714 3692
rect 31021 3689 31033 3692
rect 31067 3689 31079 3723
rect 37366 3720 37372 3732
rect 37327 3692 37372 3720
rect 31021 3683 31079 3689
rect 37366 3680 37372 3692
rect 37424 3680 37430 3732
rect 37918 3720 37924 3732
rect 37879 3692 37924 3720
rect 37918 3680 37924 3692
rect 37976 3680 37982 3732
rect 38102 3680 38108 3732
rect 38160 3720 38166 3732
rect 39577 3723 39635 3729
rect 39577 3720 39589 3723
rect 38160 3692 39589 3720
rect 38160 3680 38166 3692
rect 39577 3689 39589 3692
rect 39623 3689 39635 3723
rect 39577 3683 39635 3689
rect 19613 3655 19671 3661
rect 19613 3621 19625 3655
rect 19659 3652 19671 3655
rect 21450 3652 21456 3664
rect 19659 3624 21456 3652
rect 19659 3621 19671 3624
rect 19613 3615 19671 3621
rect 21450 3612 21456 3624
rect 21508 3612 21514 3664
rect 26970 3652 26976 3664
rect 22020 3624 26976 3652
rect 18601 3587 18659 3593
rect 18601 3553 18613 3587
rect 18647 3584 18659 3587
rect 20070 3584 20076 3596
rect 18647 3556 20076 3584
rect 18647 3553 18659 3556
rect 18601 3547 18659 3553
rect 20070 3544 20076 3556
rect 20128 3544 20134 3596
rect 22020 3593 22048 3624
rect 26970 3612 26976 3624
rect 27028 3612 27034 3664
rect 29178 3652 29184 3664
rect 28552 3624 29184 3652
rect 22005 3587 22063 3593
rect 22005 3553 22017 3587
rect 22051 3553 22063 3587
rect 22005 3547 22063 3553
rect 26053 3587 26111 3593
rect 26053 3553 26065 3587
rect 26099 3584 26111 3587
rect 28552 3584 28580 3624
rect 29178 3612 29184 3624
rect 29236 3612 29242 3664
rect 32214 3612 32220 3664
rect 32272 3652 32278 3664
rect 32272 3624 35480 3652
rect 32272 3612 32278 3624
rect 26099 3556 28580 3584
rect 28629 3587 28687 3593
rect 26099 3553 26111 3556
rect 26053 3547 26111 3553
rect 28629 3553 28641 3587
rect 28675 3584 28687 3587
rect 29638 3584 29644 3596
rect 28675 3556 29644 3584
rect 28675 3553 28687 3556
rect 28629 3547 28687 3553
rect 29638 3544 29644 3556
rect 29696 3544 29702 3596
rect 32490 3584 32496 3596
rect 32451 3556 32496 3584
rect 32490 3544 32496 3556
rect 32548 3544 32554 3596
rect 35342 3584 35348 3596
rect 34348 3556 35348 3584
rect 34348 3528 34376 3556
rect 35342 3544 35348 3556
rect 35400 3544 35406 3596
rect 35452 3593 35480 3624
rect 36630 3612 36636 3664
rect 36688 3652 36694 3664
rect 38933 3655 38991 3661
rect 38933 3652 38945 3655
rect 36688 3624 38945 3652
rect 36688 3612 36694 3624
rect 38933 3621 38945 3624
rect 38979 3621 38991 3655
rect 38933 3615 38991 3621
rect 39390 3612 39396 3664
rect 39448 3652 39454 3664
rect 40865 3655 40923 3661
rect 40865 3652 40877 3655
rect 39448 3624 40877 3652
rect 39448 3612 39454 3624
rect 40865 3621 40877 3624
rect 40911 3621 40923 3655
rect 40865 3615 40923 3621
rect 42150 3612 42156 3664
rect 42208 3652 42214 3664
rect 42889 3655 42947 3661
rect 42889 3652 42901 3655
rect 42208 3624 42901 3652
rect 42208 3612 42214 3624
rect 42889 3621 42901 3624
rect 42935 3621 42947 3655
rect 42889 3615 42947 3621
rect 43254 3612 43260 3664
rect 43312 3652 43318 3664
rect 44177 3655 44235 3661
rect 44177 3652 44189 3655
rect 43312 3624 44189 3652
rect 43312 3612 43318 3624
rect 44177 3621 44189 3624
rect 44223 3621 44235 3655
rect 44177 3615 44235 3621
rect 45462 3612 45468 3664
rect 45520 3652 45526 3664
rect 46109 3655 46167 3661
rect 46109 3652 46121 3655
rect 45520 3624 46121 3652
rect 45520 3612 45526 3624
rect 46109 3621 46121 3624
rect 46155 3621 46167 3655
rect 46109 3615 46167 3621
rect 35437 3587 35495 3593
rect 35437 3553 35449 3587
rect 35483 3553 35495 3587
rect 35437 3547 35495 3553
rect 35526 3544 35532 3596
rect 35584 3584 35590 3596
rect 35584 3556 38516 3584
rect 35584 3544 35590 3556
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 9401 3519 9459 3525
rect 9401 3516 9413 3519
rect 9364 3488 9413 3516
rect 9364 3476 9370 3488
rect 9401 3485 9413 3488
rect 9447 3485 9459 3519
rect 9401 3479 9459 3485
rect 10226 3476 10232 3528
rect 10284 3516 10290 3528
rect 10321 3519 10379 3525
rect 10321 3516 10333 3519
rect 10284 3488 10333 3516
rect 10284 3476 10290 3488
rect 10321 3485 10333 3488
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 11882 3476 11888 3528
rect 11940 3516 11946 3528
rect 11977 3519 12035 3525
rect 11977 3516 11989 3519
rect 11940 3488 11989 3516
rect 11940 3476 11946 3488
rect 11977 3485 11989 3488
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 12710 3476 12716 3528
rect 12768 3516 12774 3528
rect 12805 3519 12863 3525
rect 12805 3516 12817 3519
rect 12768 3488 12817 3516
rect 12768 3476 12774 3488
rect 12805 3485 12817 3488
rect 12851 3485 12863 3519
rect 12805 3479 12863 3485
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 13633 3519 13691 3525
rect 13633 3516 13645 3519
rect 13596 3488 13645 3516
rect 13596 3476 13602 3488
rect 13633 3485 13645 3488
rect 13679 3485 13691 3519
rect 13633 3479 13691 3485
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 14424 3488 14473 3516
rect 14424 3476 14430 3488
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 15197 3519 15255 3525
rect 15197 3516 15209 3519
rect 14976 3488 15209 3516
rect 14976 3476 14982 3488
rect 15197 3485 15209 3488
rect 15243 3485 15255 3519
rect 15197 3479 15255 3485
rect 15746 3476 15752 3528
rect 15804 3516 15810 3528
rect 15841 3519 15899 3525
rect 15841 3516 15853 3519
rect 15804 3488 15853 3516
rect 15804 3476 15810 3488
rect 15841 3485 15853 3488
rect 15887 3485 15899 3519
rect 15841 3479 15899 3485
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3516 16727 3519
rect 16850 3516 16856 3528
rect 16715 3488 16856 3516
rect 16715 3485 16727 3488
rect 16669 3479 16727 3485
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 17313 3519 17371 3525
rect 17313 3485 17325 3519
rect 17359 3516 17371 3519
rect 17862 3516 17868 3528
rect 17359 3488 17868 3516
rect 17359 3485 17371 3488
rect 17313 3479 17371 3485
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 17957 3519 18015 3525
rect 17957 3485 17969 3519
rect 18003 3516 18015 3519
rect 18138 3516 18144 3528
rect 18003 3488 18144 3516
rect 18003 3485 18015 3488
rect 17957 3479 18015 3485
rect 18138 3476 18144 3488
rect 18196 3476 18202 3528
rect 20257 3519 20315 3525
rect 20257 3485 20269 3519
rect 20303 3485 20315 3519
rect 20257 3479 20315 3485
rect 20272 3380 20300 3479
rect 22554 3476 22560 3528
rect 22612 3516 22618 3528
rect 24213 3519 24271 3525
rect 22612 3488 22657 3516
rect 22612 3476 22618 3488
rect 24213 3485 24225 3519
rect 24259 3516 24271 3519
rect 24578 3516 24584 3528
rect 24259 3488 24584 3516
rect 24259 3485 24271 3488
rect 24213 3479 24271 3485
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 26568 3488 26613 3516
rect 26568 3476 26574 3488
rect 27430 3476 27436 3528
rect 27488 3516 27494 3528
rect 27525 3519 27583 3525
rect 27525 3516 27537 3519
rect 27488 3488 27537 3516
rect 27488 3476 27494 3488
rect 27525 3485 27537 3488
rect 27571 3485 27583 3519
rect 27525 3479 27583 3485
rect 33686 3476 33692 3528
rect 33744 3516 33750 3528
rect 34330 3516 34336 3528
rect 33744 3488 33789 3516
rect 34243 3488 34336 3516
rect 33744 3476 33750 3488
rect 34330 3476 34336 3488
rect 34388 3476 34394 3528
rect 34974 3516 34980 3528
rect 34935 3488 34980 3516
rect 34974 3476 34980 3488
rect 35032 3476 35038 3528
rect 37366 3476 37372 3528
rect 37424 3516 37430 3528
rect 37461 3519 37519 3525
rect 37461 3516 37473 3519
rect 37424 3488 37473 3516
rect 37424 3476 37430 3488
rect 37461 3485 37473 3488
rect 37507 3485 37519 3519
rect 38488 3516 38516 3556
rect 38562 3544 38568 3596
rect 38620 3584 38626 3596
rect 40221 3587 40279 3593
rect 40221 3584 40233 3587
rect 38620 3556 40233 3584
rect 38620 3544 38626 3556
rect 40221 3553 40233 3556
rect 40267 3553 40279 3587
rect 40221 3547 40279 3553
rect 40770 3544 40776 3596
rect 40828 3584 40834 3596
rect 41509 3587 41567 3593
rect 41509 3584 41521 3587
rect 40828 3556 41521 3584
rect 40828 3544 40834 3556
rect 41509 3553 41521 3556
rect 41555 3553 41567 3587
rect 41509 3547 41567 3553
rect 44082 3544 44088 3596
rect 44140 3584 44146 3596
rect 44821 3587 44879 3593
rect 44821 3584 44833 3587
rect 44140 3556 44833 3584
rect 44140 3544 44146 3556
rect 44821 3553 44833 3556
rect 44867 3553 44879 3587
rect 44821 3547 44879 3553
rect 38488 3488 39528 3516
rect 37461 3479 37519 3485
rect 22373 3451 22431 3457
rect 22373 3417 22385 3451
rect 22419 3448 22431 3451
rect 23842 3448 23848 3460
rect 22419 3420 23848 3448
rect 22419 3417 22431 3420
rect 22373 3411 22431 3417
rect 23842 3408 23848 3420
rect 23900 3408 23906 3460
rect 26326 3448 26332 3460
rect 26287 3420 26332 3448
rect 26326 3408 26332 3420
rect 26384 3408 26390 3460
rect 28813 3451 28871 3457
rect 28813 3417 28825 3451
rect 28859 3448 28871 3451
rect 29086 3448 29092 3460
rect 28859 3420 29092 3448
rect 28859 3417 28871 3420
rect 28813 3411 28871 3417
rect 29086 3408 29092 3420
rect 29144 3408 29150 3460
rect 30469 3451 30527 3457
rect 30469 3417 30481 3451
rect 30515 3448 30527 3451
rect 31018 3448 31024 3460
rect 30515 3420 31024 3448
rect 30515 3417 30527 3420
rect 30469 3411 30527 3417
rect 31018 3408 31024 3420
rect 31076 3408 31082 3460
rect 33505 3451 33563 3457
rect 33505 3417 33517 3451
rect 33551 3448 33563 3451
rect 34241 3451 34299 3457
rect 34241 3448 34253 3451
rect 33551 3420 34253 3448
rect 33551 3417 33563 3420
rect 33505 3411 33563 3417
rect 34241 3417 34253 3420
rect 34287 3417 34299 3451
rect 34241 3411 34299 3417
rect 35161 3451 35219 3457
rect 35161 3417 35173 3451
rect 35207 3448 35219 3451
rect 35342 3448 35348 3460
rect 35207 3420 35348 3448
rect 35207 3417 35219 3420
rect 35161 3411 35219 3417
rect 35342 3408 35348 3420
rect 35400 3408 35406 3460
rect 36906 3408 36912 3460
rect 36964 3448 36970 3460
rect 39022 3448 39028 3460
rect 36964 3420 39028 3448
rect 36964 3408 36970 3420
rect 39022 3408 39028 3420
rect 39080 3408 39086 3460
rect 23658 3380 23664 3392
rect 20272 3352 23664 3380
rect 23658 3340 23664 3352
rect 23716 3340 23722 3392
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 38746 3380 38752 3392
rect 34848 3352 38752 3380
rect 34848 3340 34854 3352
rect 38746 3340 38752 3352
rect 38804 3340 38810 3392
rect 39500 3380 39528 3488
rect 41322 3476 41328 3528
rect 41380 3516 41386 3528
rect 42153 3519 42211 3525
rect 42153 3516 42165 3519
rect 41380 3488 42165 3516
rect 41380 3476 41386 3488
rect 42153 3485 42165 3488
rect 42199 3485 42211 3519
rect 42153 3479 42211 3485
rect 42702 3476 42708 3528
rect 42760 3516 42766 3528
rect 43533 3519 43591 3525
rect 43533 3516 43545 3519
rect 42760 3488 43545 3516
rect 42760 3476 42766 3488
rect 43533 3485 43545 3488
rect 43579 3485 43591 3519
rect 43533 3479 43591 3485
rect 44910 3476 44916 3528
rect 44968 3516 44974 3528
rect 45465 3519 45523 3525
rect 45465 3516 45477 3519
rect 44968 3488 45477 3516
rect 44968 3476 44974 3488
rect 45465 3485 45477 3488
rect 45511 3485 45523 3519
rect 45465 3479 45523 3485
rect 46290 3476 46296 3528
rect 46348 3516 46354 3528
rect 46845 3519 46903 3525
rect 46845 3516 46857 3519
rect 46348 3488 46857 3516
rect 46348 3476 46354 3488
rect 46845 3485 46857 3488
rect 46891 3485 46903 3519
rect 46845 3479 46903 3485
rect 47118 3476 47124 3528
rect 47176 3516 47182 3528
rect 47489 3519 47547 3525
rect 47489 3516 47501 3519
rect 47176 3488 47501 3516
rect 47176 3476 47182 3488
rect 47489 3485 47501 3488
rect 47535 3485 47547 3519
rect 47489 3479 47547 3485
rect 47670 3476 47676 3528
rect 47728 3516 47734 3528
rect 48133 3519 48191 3525
rect 48133 3516 48145 3519
rect 47728 3488 48145 3516
rect 47728 3476 47734 3488
rect 48133 3485 48145 3488
rect 48179 3485 48191 3519
rect 48133 3479 48191 3485
rect 49050 3476 49056 3528
rect 49108 3516 49114 3528
rect 49145 3519 49203 3525
rect 49145 3516 49157 3519
rect 49108 3488 49157 3516
rect 49108 3476 49114 3488
rect 49145 3485 49157 3488
rect 49191 3485 49203 3519
rect 49145 3479 49203 3485
rect 49602 3476 49608 3528
rect 49660 3516 49666 3528
rect 49789 3519 49847 3525
rect 49789 3516 49801 3519
rect 49660 3488 49801 3516
rect 49660 3476 49666 3488
rect 49789 3485 49801 3488
rect 49835 3485 49847 3519
rect 49789 3479 49847 3485
rect 50982 3476 50988 3528
rect 51040 3516 51046 3528
rect 51077 3519 51135 3525
rect 51077 3516 51089 3519
rect 51040 3488 51089 3516
rect 51040 3476 51046 3488
rect 51077 3485 51089 3488
rect 51123 3485 51135 3519
rect 51077 3479 51135 3485
rect 51534 3476 51540 3528
rect 51592 3516 51598 3528
rect 51721 3519 51779 3525
rect 51721 3516 51733 3519
rect 51592 3488 51733 3516
rect 51592 3476 51598 3488
rect 51721 3485 51733 3488
rect 51767 3485 51779 3519
rect 51721 3479 51779 3485
rect 40034 3380 40040 3392
rect 39500 3352 40040 3380
rect 40034 3340 40040 3352
rect 40092 3340 40098 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 21545 3179 21603 3185
rect 21545 3145 21557 3179
rect 21591 3176 21603 3179
rect 24946 3176 24952 3188
rect 21591 3148 24952 3176
rect 21591 3145 21603 3148
rect 21545 3139 21603 3145
rect 24946 3136 24952 3148
rect 25004 3136 25010 3188
rect 29454 3176 29460 3188
rect 29415 3148 29460 3176
rect 29454 3136 29460 3148
rect 29512 3136 29518 3188
rect 36354 3136 36360 3188
rect 36412 3176 36418 3188
rect 37458 3176 37464 3188
rect 36412 3148 37464 3176
rect 36412 3136 36418 3148
rect 37458 3136 37464 3148
rect 37516 3136 37522 3188
rect 19978 3068 19984 3120
rect 20036 3108 20042 3120
rect 24210 3108 24216 3120
rect 20036 3080 24216 3108
rect 20036 3068 20042 3080
rect 24210 3068 24216 3080
rect 24268 3068 24274 3120
rect 35434 3068 35440 3120
rect 35492 3108 35498 3120
rect 37185 3111 37243 3117
rect 37185 3108 37197 3111
rect 35492 3080 37197 3108
rect 35492 3068 35498 3080
rect 37185 3077 37197 3080
rect 37231 3077 37243 3111
rect 37185 3071 37243 3077
rect 37550 3068 37556 3120
rect 37608 3108 37614 3120
rect 38102 3108 38108 3120
rect 37608 3080 38108 3108
rect 37608 3068 37614 3080
rect 38102 3068 38108 3080
rect 38160 3068 38166 3120
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3040 18751 3043
rect 21174 3040 21180 3052
rect 18739 3012 21180 3040
rect 18739 3009 18751 3012
rect 18693 3003 18751 3009
rect 21174 3000 21180 3012
rect 21232 3000 21238 3052
rect 21637 3043 21695 3049
rect 21637 3009 21649 3043
rect 21683 3040 21695 3043
rect 22186 3040 22192 3052
rect 21683 3012 22192 3040
rect 21683 3009 21695 3012
rect 21637 3003 21695 3009
rect 22186 3000 22192 3012
rect 22244 3000 22250 3052
rect 22281 3043 22339 3049
rect 22281 3009 22293 3043
rect 22327 3040 22339 3043
rect 22554 3040 22560 3052
rect 22327 3012 22560 3040
rect 22327 3009 22339 3012
rect 22281 3003 22339 3009
rect 22554 3000 22560 3012
rect 22612 3000 22618 3052
rect 24578 3000 24584 3052
rect 24636 3040 24642 3052
rect 25593 3043 25651 3049
rect 24636 3012 24681 3040
rect 24636 3000 24642 3012
rect 25593 3009 25605 3043
rect 25639 3040 25651 3043
rect 26510 3040 26516 3052
rect 25639 3012 26516 3040
rect 25639 3009 25651 3012
rect 25593 3003 25651 3009
rect 26510 3000 26516 3012
rect 26568 3000 26574 3052
rect 29546 3040 29552 3052
rect 29507 3012 29552 3040
rect 29546 3000 29552 3012
rect 29604 3000 29610 3052
rect 34974 3000 34980 3052
rect 35032 3040 35038 3052
rect 35345 3043 35403 3049
rect 35345 3040 35357 3043
rect 35032 3012 35357 3040
rect 35032 3000 35038 3012
rect 35345 3009 35357 3012
rect 35391 3009 35403 3043
rect 37001 3043 37059 3049
rect 37001 3040 37013 3043
rect 35345 3003 35403 3009
rect 35866 3012 36124 3040
rect 15381 2975 15439 2981
rect 15381 2941 15393 2975
rect 15427 2972 15439 2975
rect 16022 2972 16028 2984
rect 15427 2944 16028 2972
rect 15427 2941 15439 2944
rect 15381 2935 15439 2941
rect 16022 2932 16028 2944
rect 16080 2932 16086 2984
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2972 17463 2975
rect 18966 2972 18972 2984
rect 17451 2944 18972 2972
rect 17451 2941 17463 2944
rect 17405 2935 17463 2941
rect 18966 2932 18972 2944
rect 19024 2932 19030 2984
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2972 19395 2975
rect 24121 2975 24179 2981
rect 19383 2944 22600 2972
rect 19383 2941 19395 2944
rect 19337 2935 19395 2941
rect 22572 2916 22600 2944
rect 24121 2941 24133 2975
rect 24167 2941 24179 2975
rect 24121 2935 24179 2941
rect 24397 2975 24455 2981
rect 24397 2941 24409 2975
rect 24443 2972 24455 2975
rect 25222 2972 25228 2984
rect 24443 2944 25228 2972
rect 24443 2941 24455 2944
rect 24397 2935 24455 2941
rect 18049 2907 18107 2913
rect 18049 2873 18061 2907
rect 18095 2904 18107 2907
rect 19518 2904 19524 2916
rect 18095 2876 19524 2904
rect 18095 2873 18107 2876
rect 18049 2867 18107 2873
rect 19518 2864 19524 2876
rect 19576 2864 19582 2916
rect 19978 2904 19984 2916
rect 19939 2876 19984 2904
rect 19978 2864 19984 2876
rect 20036 2864 20042 2916
rect 20625 2907 20683 2913
rect 20625 2873 20637 2907
rect 20671 2904 20683 2907
rect 20671 2876 22508 2904
rect 20671 2873 20683 2876
rect 20625 2867 20683 2873
rect 7469 2839 7527 2845
rect 7469 2805 7481 2839
rect 7515 2836 7527 2839
rect 7650 2836 7656 2848
rect 7515 2808 7656 2836
rect 7515 2805 7527 2808
rect 7469 2799 7527 2805
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 8113 2839 8171 2845
rect 8113 2805 8125 2839
rect 8159 2836 8171 2839
rect 8202 2836 8208 2848
rect 8159 2808 8208 2836
rect 8159 2805 8171 2808
rect 8113 2799 8171 2805
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 8757 2839 8815 2845
rect 8757 2805 8769 2839
rect 8803 2836 8815 2839
rect 8938 2836 8944 2848
rect 8803 2808 8944 2836
rect 8803 2805 8815 2808
rect 8757 2799 8815 2805
rect 8938 2796 8944 2808
rect 8996 2796 9002 2848
rect 9493 2839 9551 2845
rect 9493 2805 9505 2839
rect 9539 2836 9551 2839
rect 9950 2836 9956 2848
rect 9539 2808 9956 2836
rect 9539 2805 9551 2808
rect 9493 2799 9551 2805
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 10137 2839 10195 2845
rect 10137 2805 10149 2839
rect 10183 2836 10195 2839
rect 10502 2836 10508 2848
rect 10183 2808 10508 2836
rect 10183 2805 10195 2808
rect 10137 2799 10195 2805
rect 10502 2796 10508 2808
rect 10560 2796 10566 2848
rect 10781 2839 10839 2845
rect 10781 2805 10793 2839
rect 10827 2836 10839 2839
rect 11054 2836 11060 2848
rect 10827 2808 11060 2836
rect 10827 2805 10839 2808
rect 10781 2799 10839 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11425 2839 11483 2845
rect 11425 2805 11437 2839
rect 11471 2836 11483 2839
rect 11606 2836 11612 2848
rect 11471 2808 11612 2836
rect 11471 2805 11483 2808
rect 11425 2799 11483 2805
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 12069 2839 12127 2845
rect 12069 2805 12081 2839
rect 12115 2836 12127 2839
rect 12158 2836 12164 2848
rect 12115 2808 12164 2836
rect 12115 2805 12127 2808
rect 12069 2799 12127 2805
rect 12158 2796 12164 2808
rect 12216 2796 12222 2848
rect 12713 2839 12771 2845
rect 12713 2805 12725 2839
rect 12759 2836 12771 2839
rect 12986 2836 12992 2848
rect 12759 2808 12992 2836
rect 12759 2805 12771 2808
rect 12713 2799 12771 2805
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 13449 2839 13507 2845
rect 13449 2805 13461 2839
rect 13495 2836 13507 2839
rect 13814 2836 13820 2848
rect 13495 2808 13820 2836
rect 13495 2805 13507 2808
rect 13449 2799 13507 2805
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 14090 2836 14096 2848
rect 14051 2808 14096 2836
rect 14090 2796 14096 2808
rect 14148 2796 14154 2848
rect 14737 2839 14795 2845
rect 14737 2805 14749 2839
rect 14783 2836 14795 2839
rect 15194 2836 15200 2848
rect 14783 2808 15200 2836
rect 14783 2805 14795 2808
rect 14737 2799 14795 2805
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 16025 2839 16083 2845
rect 16025 2805 16037 2839
rect 16071 2836 16083 2839
rect 16574 2836 16580 2848
rect 16071 2808 16580 2836
rect 16071 2805 16083 2808
rect 16025 2799 16083 2805
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 16669 2839 16727 2845
rect 16669 2805 16681 2839
rect 16715 2836 16727 2839
rect 17310 2836 17316 2848
rect 16715 2808 17316 2836
rect 16715 2805 16727 2808
rect 16669 2799 16727 2805
rect 17310 2796 17316 2808
rect 17368 2796 17374 2848
rect 22480 2836 22508 2876
rect 22554 2864 22560 2916
rect 22612 2864 22618 2916
rect 24136 2904 24164 2935
rect 25222 2932 25228 2944
rect 25280 2932 25286 2984
rect 26237 2975 26295 2981
rect 26237 2941 26249 2975
rect 26283 2972 26295 2975
rect 26697 2975 26755 2981
rect 26697 2972 26709 2975
rect 26283 2944 26709 2972
rect 26283 2941 26295 2944
rect 26237 2935 26295 2941
rect 26697 2941 26709 2944
rect 26743 2941 26755 2975
rect 26697 2935 26755 2941
rect 26881 2975 26939 2981
rect 26881 2941 26893 2975
rect 26927 2972 26939 2975
rect 27798 2972 27804 2984
rect 26927 2944 27804 2972
rect 26927 2941 26939 2944
rect 26881 2935 26939 2941
rect 27798 2932 27804 2944
rect 27856 2932 27862 2984
rect 28537 2975 28595 2981
rect 28537 2941 28549 2975
rect 28583 2972 28595 2975
rect 29454 2972 29460 2984
rect 28583 2944 29460 2972
rect 28583 2941 28595 2944
rect 28537 2935 28595 2941
rect 29454 2932 29460 2944
rect 29512 2932 29518 2984
rect 30101 2975 30159 2981
rect 30101 2941 30113 2975
rect 30147 2941 30159 2975
rect 30101 2935 30159 2941
rect 30285 2975 30343 2981
rect 30285 2941 30297 2975
rect 30331 2972 30343 2975
rect 31110 2972 31116 2984
rect 30331 2944 31116 2972
rect 30331 2941 30343 2944
rect 30285 2935 30343 2941
rect 28902 2904 28908 2916
rect 24136 2876 28908 2904
rect 28902 2864 28908 2876
rect 28960 2864 28966 2916
rect 30116 2904 30144 2935
rect 31110 2932 31116 2944
rect 31168 2932 31174 2984
rect 31205 2975 31263 2981
rect 31205 2941 31217 2975
rect 31251 2941 31263 2975
rect 31205 2935 31263 2941
rect 30374 2904 30380 2916
rect 30116 2876 30380 2904
rect 30374 2864 30380 2876
rect 30432 2864 30438 2916
rect 30834 2864 30840 2916
rect 30892 2904 30898 2916
rect 31220 2904 31248 2935
rect 31938 2932 31944 2984
rect 31996 2972 32002 2984
rect 33045 2975 33103 2981
rect 33045 2972 33057 2975
rect 31996 2944 33057 2972
rect 31996 2932 32002 2944
rect 33045 2941 33057 2944
rect 33091 2941 33103 2975
rect 34698 2972 34704 2984
rect 34659 2944 34704 2972
rect 33045 2935 33103 2941
rect 34698 2932 34704 2944
rect 34756 2932 34762 2984
rect 34885 2975 34943 2981
rect 34885 2941 34897 2975
rect 34931 2941 34943 2975
rect 35866 2972 35894 3012
rect 34885 2935 34943 2941
rect 34992 2944 35894 2972
rect 30892 2876 31248 2904
rect 30892 2864 30898 2876
rect 34514 2864 34520 2916
rect 34572 2904 34578 2916
rect 34900 2904 34928 2935
rect 34572 2876 34928 2904
rect 34572 2864 34578 2876
rect 25038 2836 25044 2848
rect 22480 2808 25044 2836
rect 25038 2796 25044 2808
rect 25096 2796 25102 2848
rect 25406 2796 25412 2848
rect 25464 2836 25470 2848
rect 26418 2836 26424 2848
rect 25464 2808 26424 2836
rect 25464 2796 25470 2808
rect 26418 2796 26424 2808
rect 26476 2796 26482 2848
rect 33594 2796 33600 2848
rect 33652 2836 33658 2848
rect 34992 2836 35020 2944
rect 35802 2864 35808 2916
rect 35860 2904 35866 2916
rect 36096 2904 36124 3012
rect 36188 3012 37013 3040
rect 36188 2981 36216 3012
rect 37001 3009 37013 3012
rect 37047 3009 37059 3043
rect 37001 3003 37059 3009
rect 38378 3000 38384 3052
rect 38436 3040 38442 3052
rect 40957 3043 41015 3049
rect 40957 3040 40969 3043
rect 38436 3012 40969 3040
rect 38436 3000 38442 3012
rect 40957 3009 40969 3012
rect 41003 3009 41015 3043
rect 40957 3003 41015 3009
rect 41046 3000 41052 3052
rect 41104 3040 41110 3052
rect 42889 3043 42947 3049
rect 42889 3040 42901 3043
rect 41104 3012 42901 3040
rect 41104 3000 41110 3012
rect 42889 3009 42901 3012
rect 42935 3009 42947 3043
rect 42889 3003 42947 3009
rect 36173 2975 36231 2981
rect 36173 2941 36185 2975
rect 36219 2941 36231 2975
rect 36173 2935 36231 2941
rect 37645 2975 37703 2981
rect 37645 2941 37657 2975
rect 37691 2941 37703 2975
rect 37645 2935 37703 2941
rect 37660 2904 37688 2935
rect 39666 2932 39672 2984
rect 39724 2972 39730 2984
rect 41601 2975 41659 2981
rect 41601 2972 41613 2975
rect 39724 2944 41613 2972
rect 39724 2932 39730 2944
rect 41601 2941 41613 2944
rect 41647 2941 41659 2975
rect 41601 2935 41659 2941
rect 41874 2932 41880 2984
rect 41932 2972 41938 2984
rect 43533 2975 43591 2981
rect 43533 2972 43545 2975
rect 41932 2944 43545 2972
rect 41932 2932 41938 2944
rect 43533 2941 43545 2944
rect 43579 2941 43591 2975
rect 43533 2935 43591 2941
rect 44358 2932 44364 2984
rect 44416 2972 44422 2984
rect 45557 2975 45615 2981
rect 45557 2972 45569 2975
rect 44416 2944 45569 2972
rect 44416 2932 44422 2944
rect 45557 2941 45569 2944
rect 45603 2941 45615 2975
rect 45557 2935 45615 2941
rect 46566 2932 46572 2984
rect 46624 2972 46630 2984
rect 47489 2975 47547 2981
rect 47489 2972 47501 2975
rect 46624 2944 47501 2972
rect 46624 2932 46630 2944
rect 47489 2941 47501 2944
rect 47535 2941 47547 2975
rect 47489 2935 47547 2941
rect 49878 2932 49884 2984
rect 49936 2972 49942 2984
rect 50801 2975 50859 2981
rect 50801 2972 50813 2975
rect 49936 2944 50813 2972
rect 49936 2932 49942 2944
rect 50801 2941 50813 2944
rect 50847 2941 50859 2975
rect 50801 2935 50859 2941
rect 52086 2932 52092 2984
rect 52144 2972 52150 2984
rect 52825 2975 52883 2981
rect 52825 2972 52837 2975
rect 52144 2944 52837 2972
rect 52144 2932 52150 2944
rect 52825 2941 52837 2944
rect 52871 2941 52883 2975
rect 52825 2935 52883 2941
rect 35860 2876 36032 2904
rect 36096 2876 37688 2904
rect 35860 2864 35866 2876
rect 33652 2808 35020 2836
rect 33652 2796 33658 2808
rect 35434 2796 35440 2848
rect 35492 2836 35498 2848
rect 35894 2836 35900 2848
rect 35492 2808 35900 2836
rect 35492 2796 35498 2808
rect 35894 2796 35900 2808
rect 35952 2796 35958 2848
rect 36004 2836 36032 2876
rect 38010 2864 38016 2916
rect 38068 2904 38074 2916
rect 38930 2904 38936 2916
rect 38068 2876 38936 2904
rect 38068 2864 38074 2876
rect 38930 2864 38936 2876
rect 38988 2864 38994 2916
rect 39022 2864 39028 2916
rect 39080 2904 39086 2916
rect 39945 2907 40003 2913
rect 39945 2904 39957 2907
rect 39080 2876 39957 2904
rect 39080 2864 39086 2876
rect 39945 2873 39957 2876
rect 39991 2873 40003 2907
rect 39945 2867 40003 2873
rect 40494 2864 40500 2916
rect 40552 2904 40558 2916
rect 42245 2907 42303 2913
rect 42245 2904 42257 2907
rect 40552 2876 42257 2904
rect 40552 2864 40558 2876
rect 42245 2873 42257 2876
rect 42291 2873 42303 2907
rect 42245 2867 42303 2873
rect 42978 2864 42984 2916
rect 43036 2904 43042 2916
rect 44177 2907 44235 2913
rect 44177 2904 44189 2907
rect 43036 2876 44189 2904
rect 43036 2864 43042 2876
rect 44177 2873 44189 2876
rect 44223 2873 44235 2907
rect 44177 2867 44235 2873
rect 45186 2864 45192 2916
rect 45244 2904 45250 2916
rect 46201 2907 46259 2913
rect 46201 2904 46213 2907
rect 45244 2876 46213 2904
rect 45244 2864 45250 2876
rect 46201 2873 46213 2876
rect 46247 2873 46259 2907
rect 46201 2867 46259 2873
rect 47394 2864 47400 2916
rect 47452 2904 47458 2916
rect 48133 2907 48191 2913
rect 48133 2904 48145 2907
rect 47452 2876 48145 2904
rect 47452 2864 47458 2876
rect 48133 2873 48145 2876
rect 48179 2873 48191 2907
rect 48133 2867 48191 2873
rect 48774 2864 48780 2916
rect 48832 2904 48838 2916
rect 49513 2907 49571 2913
rect 49513 2904 49525 2907
rect 48832 2876 49525 2904
rect 48832 2864 48838 2876
rect 49513 2873 49525 2876
rect 49559 2873 49571 2907
rect 49513 2867 49571 2873
rect 50706 2864 50712 2916
rect 50764 2904 50770 2916
rect 51445 2907 51503 2913
rect 51445 2904 51457 2907
rect 50764 2876 51457 2904
rect 50764 2864 50770 2876
rect 51445 2873 51457 2876
rect 51491 2873 51503 2907
rect 51445 2867 51503 2873
rect 39301 2839 39359 2845
rect 39301 2836 39313 2839
rect 36004 2808 39313 2836
rect 39301 2805 39313 2808
rect 39347 2805 39359 2839
rect 39301 2799 39359 2805
rect 43622 2796 43628 2848
rect 43680 2836 43686 2848
rect 44913 2839 44971 2845
rect 44913 2836 44925 2839
rect 43680 2808 44925 2836
rect 43680 2796 43686 2808
rect 44913 2805 44925 2808
rect 44959 2805 44971 2839
rect 44913 2799 44971 2805
rect 45738 2796 45744 2848
rect 45796 2836 45802 2848
rect 46845 2839 46903 2845
rect 46845 2836 46857 2839
rect 45796 2808 46857 2836
rect 45796 2796 45802 2808
rect 46845 2805 46857 2808
rect 46891 2805 46903 2839
rect 46845 2799 46903 2805
rect 47946 2796 47952 2848
rect 48004 2836 48010 2848
rect 48869 2839 48927 2845
rect 48869 2836 48881 2839
rect 48004 2808 48881 2836
rect 48004 2796 48010 2808
rect 48869 2805 48881 2808
rect 48915 2805 48927 2839
rect 48869 2799 48927 2805
rect 49326 2796 49332 2848
rect 49384 2836 49390 2848
rect 50157 2839 50215 2845
rect 50157 2836 50169 2839
rect 49384 2808 50169 2836
rect 49384 2796 49390 2808
rect 50157 2805 50169 2808
rect 50203 2805 50215 2839
rect 50157 2799 50215 2805
rect 51258 2796 51264 2848
rect 51316 2836 51322 2848
rect 52089 2839 52147 2845
rect 52089 2836 52101 2839
rect 51316 2808 52101 2836
rect 51316 2796 51322 2808
rect 52089 2805 52101 2808
rect 52135 2805 52147 2839
rect 52089 2799 52147 2805
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 22922 2592 22928 2644
rect 22980 2632 22986 2644
rect 23293 2635 23351 2641
rect 23293 2632 23305 2635
rect 22980 2604 23305 2632
rect 22980 2592 22986 2604
rect 23293 2601 23305 2604
rect 23339 2601 23351 2635
rect 23293 2595 23351 2601
rect 23842 2592 23848 2644
rect 23900 2632 23906 2644
rect 23937 2635 23995 2641
rect 23937 2632 23949 2635
rect 23900 2604 23949 2632
rect 23900 2592 23906 2604
rect 23937 2601 23949 2604
rect 23983 2601 23995 2635
rect 25222 2632 25228 2644
rect 25183 2604 25228 2632
rect 23937 2595 23995 2601
rect 25222 2592 25228 2604
rect 25280 2592 25286 2644
rect 26326 2592 26332 2644
rect 26384 2632 26390 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 26384 2604 27169 2632
rect 26384 2592 26390 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 27798 2632 27804 2644
rect 27759 2604 27804 2632
rect 27157 2595 27215 2601
rect 27798 2592 27804 2604
rect 27856 2592 27862 2644
rect 29086 2632 29092 2644
rect 29047 2604 29092 2632
rect 29086 2592 29092 2604
rect 29144 2592 29150 2644
rect 29638 2632 29644 2644
rect 29599 2604 29644 2632
rect 29638 2592 29644 2604
rect 29696 2592 29702 2644
rect 30374 2632 30380 2644
rect 30335 2604 30380 2632
rect 30374 2592 30380 2604
rect 30432 2592 30438 2644
rect 31110 2632 31116 2644
rect 31071 2604 31116 2632
rect 31110 2592 31116 2604
rect 31168 2592 31174 2644
rect 32493 2635 32551 2641
rect 32493 2601 32505 2635
rect 32539 2632 32551 2635
rect 33686 2632 33692 2644
rect 32539 2604 33692 2632
rect 32539 2601 32551 2604
rect 32493 2595 32551 2601
rect 33686 2592 33692 2604
rect 33744 2592 33750 2644
rect 34333 2635 34391 2641
rect 34333 2601 34345 2635
rect 34379 2632 34391 2635
rect 34698 2632 34704 2644
rect 34379 2604 34704 2632
rect 34379 2601 34391 2604
rect 34333 2595 34391 2601
rect 34698 2592 34704 2604
rect 34756 2592 34762 2644
rect 34977 2635 35035 2641
rect 34977 2601 34989 2635
rect 35023 2632 35035 2635
rect 35342 2632 35348 2644
rect 35023 2604 35348 2632
rect 35023 2601 35035 2604
rect 34977 2595 35035 2601
rect 35342 2592 35348 2604
rect 35400 2592 35406 2644
rect 36357 2635 36415 2641
rect 36357 2601 36369 2635
rect 36403 2632 36415 2635
rect 36998 2632 37004 2644
rect 36403 2604 37004 2632
rect 36403 2601 36415 2604
rect 36357 2595 36415 2601
rect 36998 2592 37004 2604
rect 37056 2592 37062 2644
rect 38194 2632 38200 2644
rect 38155 2604 38200 2632
rect 38194 2592 38200 2604
rect 38252 2592 38258 2644
rect 38746 2632 38752 2644
rect 38707 2604 38752 2632
rect 38746 2592 38752 2604
rect 38804 2592 38810 2644
rect 40034 2632 40040 2644
rect 39995 2604 40040 2632
rect 40034 2592 40040 2604
rect 40092 2592 40098 2644
rect 7929 2567 7987 2573
rect 7929 2533 7941 2567
rect 7975 2564 7987 2567
rect 8570 2564 8576 2576
rect 7975 2536 8576 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 8570 2524 8576 2536
rect 8628 2524 8634 2576
rect 11793 2567 11851 2573
rect 11793 2533 11805 2567
rect 11839 2564 11851 2567
rect 12434 2564 12440 2576
rect 11839 2536 12440 2564
rect 11839 2533 11851 2536
rect 11793 2527 11851 2533
rect 12434 2524 12440 2536
rect 12492 2524 12498 2576
rect 16301 2567 16359 2573
rect 16301 2533 16313 2567
rect 16347 2564 16359 2567
rect 18690 2564 18696 2576
rect 16347 2536 18696 2564
rect 16347 2533 16359 2536
rect 16301 2527 16359 2533
rect 18690 2524 18696 2536
rect 18748 2524 18754 2576
rect 21453 2567 21511 2573
rect 21453 2533 21465 2567
rect 21499 2564 21511 2567
rect 25590 2564 25596 2576
rect 21499 2536 25596 2564
rect 21499 2533 21511 2536
rect 21453 2527 21511 2533
rect 25590 2524 25596 2536
rect 25648 2524 25654 2576
rect 33137 2567 33195 2573
rect 33137 2533 33149 2567
rect 33183 2564 33195 2567
rect 34514 2564 34520 2576
rect 33183 2536 34520 2564
rect 33183 2533 33195 2536
rect 33137 2527 33195 2533
rect 34514 2524 34520 2536
rect 34572 2524 34578 2576
rect 36909 2567 36967 2573
rect 36909 2533 36921 2567
rect 36955 2564 36967 2567
rect 37182 2564 37188 2576
rect 36955 2536 37188 2564
rect 36955 2533 36967 2536
rect 36909 2527 36967 2533
rect 37182 2524 37188 2536
rect 37240 2524 37246 2576
rect 39942 2524 39948 2576
rect 40000 2564 40006 2576
rect 42613 2567 42671 2573
rect 42613 2564 42625 2567
rect 40000 2536 42625 2564
rect 40000 2524 40006 2536
rect 42613 2533 42625 2536
rect 42659 2533 42671 2567
rect 42613 2527 42671 2533
rect 43806 2524 43812 2576
rect 43864 2564 43870 2576
rect 45833 2567 45891 2573
rect 45833 2564 45845 2567
rect 43864 2536 45845 2564
rect 43864 2524 43870 2536
rect 45833 2533 45845 2536
rect 45879 2533 45891 2567
rect 45833 2527 45891 2533
rect 46842 2524 46848 2576
rect 46900 2564 46906 2576
rect 48409 2567 48467 2573
rect 48409 2564 48421 2567
rect 46900 2536 48421 2564
rect 46900 2524 46906 2536
rect 48409 2533 48421 2536
rect 48455 2533 48467 2567
rect 48409 2527 48467 2533
rect 51810 2524 51816 2576
rect 51868 2564 51874 2576
rect 53561 2567 53619 2573
rect 53561 2564 53573 2567
rect 51868 2536 53573 2564
rect 51868 2524 51874 2536
rect 53561 2533 53573 2536
rect 53607 2533 53619 2567
rect 53561 2527 53619 2533
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2496 9919 2499
rect 10778 2496 10784 2508
rect 9907 2468 10784 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2496 13783 2499
rect 14642 2496 14648 2508
rect 13771 2468 14648 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 14642 2456 14648 2468
rect 14700 2456 14706 2508
rect 15657 2499 15715 2505
rect 15657 2465 15669 2499
rect 15703 2496 15715 2499
rect 17126 2496 17132 2508
rect 15703 2468 17132 2496
rect 15703 2465 15715 2468
rect 15657 2459 15715 2465
rect 17126 2456 17132 2468
rect 17184 2456 17190 2508
rect 17589 2499 17647 2505
rect 17589 2465 17601 2499
rect 17635 2496 17647 2499
rect 20898 2496 20904 2508
rect 17635 2468 20904 2496
rect 17635 2465 17647 2468
rect 17589 2459 17647 2465
rect 20898 2456 20904 2468
rect 20956 2456 20962 2508
rect 22097 2499 22155 2505
rect 22097 2465 22109 2499
rect 22143 2496 22155 2499
rect 25866 2496 25872 2508
rect 22143 2468 25872 2496
rect 22143 2465 22155 2468
rect 22097 2459 22155 2465
rect 25866 2456 25872 2468
rect 25924 2456 25930 2508
rect 38838 2456 38844 2508
rect 38896 2496 38902 2508
rect 41969 2499 42027 2505
rect 41969 2496 41981 2499
rect 38896 2468 41981 2496
rect 38896 2456 38902 2468
rect 41969 2465 41981 2468
rect 42015 2465 42027 2499
rect 41969 2459 42027 2465
rect 42426 2456 42432 2508
rect 42484 2496 42490 2508
rect 44545 2499 44603 2505
rect 44545 2496 44557 2499
rect 42484 2468 44557 2496
rect 42484 2456 42490 2468
rect 44545 2465 44557 2468
rect 44591 2465 44603 2499
rect 44545 2459 44603 2465
rect 44634 2456 44640 2508
rect 44692 2496 44698 2508
rect 46477 2499 46535 2505
rect 46477 2496 46489 2499
rect 44692 2468 46489 2496
rect 44692 2456 44698 2468
rect 46477 2465 46489 2468
rect 46523 2465 46535 2499
rect 46477 2459 46535 2465
rect 48222 2456 48228 2508
rect 48280 2496 48286 2508
rect 49697 2499 49755 2505
rect 49697 2496 49709 2499
rect 48280 2468 49709 2496
rect 48280 2456 48286 2468
rect 49697 2465 49709 2468
rect 49743 2465 49755 2499
rect 49697 2459 49755 2465
rect 50154 2456 50160 2508
rect 50212 2496 50218 2508
rect 51629 2499 51687 2505
rect 51629 2496 51641 2499
rect 50212 2468 51641 2496
rect 50212 2456 50218 2468
rect 51629 2465 51641 2468
rect 51675 2465 51687 2499
rect 51629 2459 51687 2465
rect 52362 2456 52368 2508
rect 52420 2496 52426 2508
rect 54205 2499 54263 2505
rect 54205 2496 54217 2499
rect 52420 2468 54217 2496
rect 52420 2456 52426 2468
rect 54205 2465 54217 2468
rect 54251 2465 54263 2499
rect 54205 2459 54263 2465
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 9674 2428 9680 2440
rect 8619 2400 9680 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 11330 2428 11336 2440
rect 10551 2400 11336 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 11330 2388 11336 2400
rect 11388 2388 11394 2440
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 13262 2428 13268 2440
rect 12483 2400 13268 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2428 14427 2431
rect 15470 2428 15476 2440
rect 14415 2400 15476 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2397 18291 2431
rect 18233 2391 18291 2397
rect 19521 2431 19579 2437
rect 19521 2397 19533 2431
rect 19567 2428 19579 2431
rect 19978 2428 19984 2440
rect 19567 2400 19984 2428
rect 19567 2397 19579 2400
rect 19521 2391 19579 2397
rect 18248 2360 18276 2391
rect 19978 2388 19984 2400
rect 20036 2388 20042 2440
rect 20165 2431 20223 2437
rect 20165 2397 20177 2431
rect 20211 2428 20223 2431
rect 23290 2428 23296 2440
rect 20211 2400 23296 2428
rect 20211 2397 20223 2400
rect 20165 2391 20223 2397
rect 23290 2388 23296 2400
rect 23348 2388 23354 2440
rect 23385 2431 23443 2437
rect 23385 2397 23397 2431
rect 23431 2428 23443 2431
rect 24029 2431 24087 2437
rect 24029 2428 24041 2431
rect 23431 2400 24041 2428
rect 23431 2397 23443 2400
rect 23385 2391 23443 2397
rect 24029 2397 24041 2400
rect 24075 2428 24087 2431
rect 25317 2431 25375 2437
rect 25317 2428 25329 2431
rect 24075 2400 25329 2428
rect 24075 2397 24087 2400
rect 24029 2391 24087 2397
rect 25317 2397 25329 2400
rect 25363 2428 25375 2431
rect 25777 2431 25835 2437
rect 25777 2428 25789 2431
rect 25363 2400 25789 2428
rect 25363 2397 25375 2400
rect 25317 2391 25375 2397
rect 25777 2397 25789 2400
rect 25823 2397 25835 2431
rect 25777 2391 25835 2397
rect 27249 2431 27307 2437
rect 27249 2397 27261 2431
rect 27295 2428 27307 2431
rect 27430 2428 27436 2440
rect 27295 2400 27436 2428
rect 27295 2397 27307 2400
rect 27249 2391 27307 2397
rect 22278 2360 22284 2372
rect 18248 2332 22284 2360
rect 22278 2320 22284 2332
rect 22336 2320 22342 2372
rect 23400 2360 23428 2391
rect 27430 2388 27436 2400
rect 27488 2428 27494 2440
rect 27893 2431 27951 2437
rect 27893 2428 27905 2431
rect 27488 2400 27905 2428
rect 27488 2388 27494 2400
rect 27893 2397 27905 2400
rect 27939 2428 27951 2431
rect 29181 2431 29239 2437
rect 29181 2428 29193 2431
rect 27939 2400 29193 2428
rect 27939 2397 27951 2400
rect 27893 2391 27951 2397
rect 29181 2397 29193 2400
rect 29227 2428 29239 2431
rect 29546 2428 29552 2440
rect 29227 2400 29552 2428
rect 29227 2397 29239 2400
rect 29181 2391 29239 2397
rect 29546 2388 29552 2400
rect 29604 2428 29610 2440
rect 31205 2431 31263 2437
rect 31205 2428 31217 2431
rect 29604 2400 31217 2428
rect 29604 2388 29610 2400
rect 31205 2397 31217 2400
rect 31251 2397 31263 2431
rect 31205 2391 31263 2397
rect 34330 2388 34336 2440
rect 34388 2428 34394 2440
rect 34425 2431 34483 2437
rect 34425 2428 34437 2431
rect 34388 2400 34437 2428
rect 34388 2388 34394 2400
rect 34425 2397 34437 2400
rect 34471 2428 34483 2431
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34471 2400 34897 2428
rect 34471 2397 34483 2400
rect 34425 2391 34483 2397
rect 34885 2397 34897 2400
rect 34931 2428 34943 2431
rect 36817 2431 36875 2437
rect 36817 2428 36829 2431
rect 34931 2400 36829 2428
rect 34931 2397 34943 2400
rect 34885 2391 34943 2397
rect 36817 2397 36829 2400
rect 36863 2428 36875 2431
rect 37366 2428 37372 2440
rect 36863 2400 37372 2428
rect 36863 2397 36875 2400
rect 36817 2391 36875 2397
rect 37366 2388 37372 2400
rect 37424 2428 37430 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 37424 2400 38117 2428
rect 37424 2388 37430 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 40681 2431 40739 2437
rect 40681 2397 40693 2431
rect 40727 2397 40739 2431
rect 40681 2391 40739 2397
rect 43901 2431 43959 2437
rect 43901 2397 43913 2431
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 23216 2332 23428 2360
rect 25869 2363 25927 2369
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19518 2292 19524 2304
rect 19392 2264 19524 2292
rect 19392 2252 19398 2264
rect 19518 2252 19524 2264
rect 19576 2252 19582 2304
rect 22186 2252 22192 2304
rect 22244 2292 22250 2304
rect 23216 2292 23244 2332
rect 25869 2329 25881 2363
rect 25915 2360 25927 2363
rect 28166 2360 28172 2372
rect 25915 2332 28172 2360
rect 25915 2329 25927 2332
rect 25869 2323 25927 2329
rect 28166 2320 28172 2332
rect 28224 2320 28230 2372
rect 36078 2320 36084 2372
rect 36136 2360 36142 2372
rect 40696 2360 40724 2391
rect 36136 2332 40724 2360
rect 36136 2320 36142 2332
rect 41598 2320 41604 2372
rect 41656 2360 41662 2372
rect 43916 2360 43944 2391
rect 46014 2388 46020 2440
rect 46072 2428 46078 2440
rect 47765 2431 47823 2437
rect 47765 2428 47777 2431
rect 46072 2400 47777 2428
rect 46072 2388 46078 2400
rect 47765 2397 47777 2400
rect 47811 2397 47823 2431
rect 47765 2391 47823 2397
rect 48498 2388 48504 2440
rect 48556 2428 48562 2440
rect 50341 2431 50399 2437
rect 50341 2428 50353 2431
rect 48556 2400 50353 2428
rect 48556 2388 48562 2400
rect 50341 2397 50353 2400
rect 50387 2397 50399 2431
rect 50341 2391 50399 2397
rect 50614 2388 50620 2440
rect 50672 2428 50678 2440
rect 52273 2431 52331 2437
rect 52273 2428 52285 2431
rect 50672 2400 52285 2428
rect 50672 2388 50678 2400
rect 52273 2397 52285 2400
rect 52319 2397 52331 2431
rect 52273 2391 52331 2397
rect 41656 2332 43944 2360
rect 41656 2320 41662 2332
rect 22244 2264 23244 2292
rect 22244 2252 22250 2264
rect 23290 2252 23296 2304
rect 23348 2292 23354 2304
rect 25314 2292 25320 2304
rect 23348 2264 25320 2292
rect 23348 2252 23354 2264
rect 25314 2252 25320 2264
rect 25372 2252 25378 2304
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 19978 2048 19984 2100
rect 20036 2088 20042 2100
rect 24762 2088 24768 2100
rect 20036 2060 24768 2088
rect 20036 2048 20042 2060
rect 24762 2048 24768 2060
rect 24820 2048 24826 2100
<< via1 >>
rect 15200 57876 15252 57928
rect 25688 57876 25740 57928
rect 27620 57876 27672 57928
rect 35992 57876 36044 57928
rect 22008 57808 22060 57860
rect 24676 57808 24728 57860
rect 24768 57808 24820 57860
rect 40040 57808 40092 57860
rect 40132 57808 40184 57860
rect 20996 57740 21048 57792
rect 25044 57740 25096 57792
rect 27988 57740 28040 57792
rect 35532 57740 35584 57792
rect 35716 57740 35768 57792
rect 40408 57740 40460 57792
rect 42340 57808 42392 57860
rect 44732 57808 44784 57860
rect 49148 57740 49200 57792
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 5080 57536 5132 57588
rect 11060 57536 11112 57588
rect 11980 57536 12032 57588
rect 13360 57536 13412 57588
rect 14740 57536 14792 57588
rect 16120 57536 16172 57588
rect 17500 57536 17552 57588
rect 18880 57536 18932 57588
rect 20260 57536 20312 57588
rect 21640 57536 21692 57588
rect 23020 57536 23072 57588
rect 24400 57536 24452 57588
rect 24676 57536 24728 57588
rect 25964 57536 26016 57588
rect 27068 57536 27120 57588
rect 31300 57536 31352 57588
rect 34244 57536 34296 57588
rect 40040 57579 40092 57588
rect 40040 57545 40049 57579
rect 40049 57545 40083 57579
rect 40083 57545 40092 57579
rect 40040 57536 40092 57545
rect 3700 57468 3752 57520
rect 4620 57400 4672 57452
rect 6460 57443 6512 57452
rect 6460 57409 6469 57443
rect 6469 57409 6503 57443
rect 6503 57409 6512 57443
rect 6460 57400 6512 57409
rect 7840 57400 7892 57452
rect 8760 57400 8812 57452
rect 9220 57400 9272 57452
rect 10140 57400 10192 57452
rect 11336 57443 11388 57452
rect 11336 57409 11345 57443
rect 11345 57409 11379 57443
rect 11379 57409 11388 57443
rect 11336 57400 11388 57409
rect 12348 57443 12400 57452
rect 12348 57409 12357 57443
rect 12357 57409 12391 57443
rect 12391 57409 12400 57443
rect 12348 57400 12400 57409
rect 23204 57468 23256 57520
rect 14280 57400 14332 57452
rect 15200 57443 15252 57452
rect 15200 57409 15209 57443
rect 15209 57409 15243 57443
rect 15243 57409 15252 57443
rect 15200 57400 15252 57409
rect 15660 57400 15712 57452
rect 19248 57443 19300 57452
rect 7288 57332 7340 57384
rect 16948 57264 17000 57316
rect 7288 57239 7340 57248
rect 7288 57205 7297 57239
rect 7297 57205 7331 57239
rect 7331 57205 7340 57239
rect 7288 57196 7340 57205
rect 19248 57409 19257 57443
rect 19257 57409 19291 57443
rect 19291 57409 19300 57443
rect 19248 57400 19300 57409
rect 19984 57400 20036 57452
rect 20996 57443 21048 57452
rect 20996 57409 21005 57443
rect 21005 57409 21039 57443
rect 21039 57409 21048 57443
rect 20996 57400 21048 57409
rect 22008 57443 22060 57452
rect 22008 57409 22017 57443
rect 22017 57409 22051 57443
rect 22051 57409 22060 57443
rect 22008 57400 22060 57409
rect 23756 57443 23808 57452
rect 23756 57409 23765 57443
rect 23765 57409 23799 57443
rect 23799 57409 23808 57443
rect 23756 57400 23808 57409
rect 24768 57443 24820 57452
rect 24768 57409 24777 57443
rect 24777 57409 24811 57443
rect 24811 57409 24820 57443
rect 24768 57400 24820 57409
rect 25596 57443 25648 57452
rect 25596 57409 25605 57443
rect 25605 57409 25639 57443
rect 25639 57409 25648 57443
rect 25596 57400 25648 57409
rect 26424 57400 26476 57452
rect 27620 57443 27672 57452
rect 27620 57409 27629 57443
rect 27629 57409 27663 57443
rect 27663 57409 27672 57443
rect 27620 57400 27672 57409
rect 27896 57443 27948 57452
rect 27896 57409 27905 57443
rect 27905 57409 27939 57443
rect 27939 57409 27948 57443
rect 27896 57400 27948 57409
rect 29184 57400 29236 57452
rect 29276 57443 29328 57452
rect 29276 57409 29285 57443
rect 29285 57409 29319 57443
rect 29319 57409 29328 57443
rect 29276 57400 29328 57409
rect 33692 57468 33744 57520
rect 34520 57468 34572 57520
rect 43352 57536 43404 57588
rect 40408 57468 40460 57520
rect 52460 57468 52512 57520
rect 52828 57468 52880 57520
rect 31392 57443 31444 57452
rect 21364 57264 21416 57316
rect 26148 57332 26200 57384
rect 22468 57196 22520 57248
rect 22652 57196 22704 57248
rect 28264 57264 28316 57316
rect 28540 57332 28592 57384
rect 30012 57332 30064 57384
rect 31392 57409 31401 57443
rect 31401 57409 31435 57443
rect 31435 57409 31444 57443
rect 31392 57400 31444 57409
rect 31760 57400 31812 57452
rect 37556 57400 37608 57452
rect 40132 57400 40184 57452
rect 40868 57400 40920 57452
rect 41236 57443 41288 57452
rect 41236 57409 41245 57443
rect 41245 57409 41279 57443
rect 41279 57409 41288 57443
rect 41236 57400 41288 57409
rect 41328 57400 41380 57452
rect 31668 57375 31720 57384
rect 31668 57341 31677 57375
rect 31677 57341 31711 57375
rect 31711 57341 31720 57375
rect 31668 57332 31720 57341
rect 32588 57375 32640 57384
rect 32588 57341 32597 57375
rect 32597 57341 32631 57375
rect 32631 57341 32640 57375
rect 32588 57332 32640 57341
rect 33140 57332 33192 57384
rect 35808 57332 35860 57384
rect 35900 57332 35952 57384
rect 36176 57375 36228 57384
rect 36176 57341 36185 57375
rect 36185 57341 36219 57375
rect 36219 57341 36228 57375
rect 36176 57332 36228 57341
rect 25228 57196 25280 57248
rect 25504 57196 25556 57248
rect 27712 57239 27764 57248
rect 27712 57205 27721 57239
rect 27721 57205 27755 57239
rect 27755 57205 27764 57239
rect 27712 57196 27764 57205
rect 28356 57196 28408 57248
rect 34428 57264 34480 57316
rect 37280 57332 37332 57384
rect 38292 57332 38344 57384
rect 31208 57239 31260 57248
rect 31208 57205 31217 57239
rect 31217 57205 31251 57239
rect 31251 57205 31260 57239
rect 31208 57196 31260 57205
rect 32036 57196 32088 57248
rect 33876 57196 33928 57248
rect 34612 57196 34664 57248
rect 35348 57239 35400 57248
rect 35348 57205 35357 57239
rect 35357 57205 35391 57239
rect 35391 57205 35400 57239
rect 35348 57196 35400 57205
rect 37280 57196 37332 57248
rect 39948 57332 40000 57384
rect 40500 57375 40552 57384
rect 40500 57341 40509 57375
rect 40509 57341 40543 57375
rect 40543 57341 40552 57375
rect 42800 57400 42852 57452
rect 43536 57400 43588 57452
rect 44916 57400 44968 57452
rect 45560 57400 45612 57452
rect 46388 57400 46440 57452
rect 46756 57443 46808 57452
rect 46756 57409 46765 57443
rect 46765 57409 46799 57443
rect 46799 57409 46808 57443
rect 46756 57400 46808 57409
rect 46940 57400 46992 57452
rect 47584 57400 47636 57452
rect 49700 57400 49752 57452
rect 51080 57400 51132 57452
rect 51448 57400 51500 57452
rect 53840 57400 53892 57452
rect 54300 57400 54352 57452
rect 55220 57400 55272 57452
rect 55680 57400 55732 57452
rect 40500 57332 40552 57341
rect 43996 57332 44048 57384
rect 44456 57332 44508 57384
rect 40960 57264 41012 57316
rect 43168 57264 43220 57316
rect 40132 57196 40184 57248
rect 43904 57239 43956 57248
rect 43904 57205 43913 57239
rect 43913 57205 43947 57239
rect 43947 57205 43956 57239
rect 43904 57196 43956 57205
rect 44272 57239 44324 57248
rect 44272 57205 44281 57239
rect 44281 57205 44315 57239
rect 44315 57205 44324 57239
rect 44272 57196 44324 57205
rect 44824 57239 44876 57248
rect 44824 57205 44833 57239
rect 44833 57205 44867 57239
rect 44867 57205 44876 57239
rect 44824 57196 44876 57205
rect 45928 57239 45980 57248
rect 45928 57205 45937 57239
rect 45937 57205 45971 57239
rect 45971 57205 45980 57239
rect 45928 57196 45980 57205
rect 46388 57264 46440 57316
rect 49148 57264 49200 57316
rect 54116 57239 54168 57248
rect 54116 57205 54125 57239
rect 54125 57205 54159 57239
rect 54159 57205 54168 57239
rect 54116 57196 54168 57205
rect 54208 57196 54260 57248
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 3700 57035 3752 57044
rect 3700 57001 3709 57035
rect 3709 57001 3743 57035
rect 3743 57001 3752 57035
rect 3700 56992 3752 57001
rect 6000 56992 6052 57044
rect 7380 56992 7432 57044
rect 11520 56992 11572 57044
rect 12900 56992 12952 57044
rect 17040 56992 17092 57044
rect 18420 56992 18472 57044
rect 21180 56992 21232 57044
rect 23204 56992 23256 57044
rect 25688 57035 25740 57044
rect 25688 57001 25697 57035
rect 25697 57001 25731 57035
rect 25731 57001 25740 57035
rect 25688 56992 25740 57001
rect 26976 56992 27028 57044
rect 29828 56992 29880 57044
rect 30012 56992 30064 57044
rect 30840 56992 30892 57044
rect 31392 56992 31444 57044
rect 34244 57035 34296 57044
rect 34244 57001 34253 57035
rect 34253 57001 34287 57035
rect 34287 57001 34296 57035
rect 34244 56992 34296 57001
rect 34704 56992 34756 57044
rect 36728 56992 36780 57044
rect 39856 56992 39908 57044
rect 41788 56992 41840 57044
rect 44272 56992 44324 57044
rect 46020 56992 46072 57044
rect 47860 56992 47912 57044
rect 50160 56992 50212 57044
rect 51540 56992 51592 57044
rect 52460 56992 52512 57044
rect 52920 56992 52972 57044
rect 53472 56992 53524 57044
rect 54760 56992 54812 57044
rect 55220 56992 55272 57044
rect 56140 56992 56192 57044
rect 19248 56924 19300 56976
rect 11336 56856 11388 56908
rect 21364 56856 21416 56908
rect 22468 56924 22520 56976
rect 30288 56924 30340 56976
rect 24032 56856 24084 56908
rect 24860 56856 24912 56908
rect 25044 56899 25096 56908
rect 25044 56865 25053 56899
rect 25053 56865 25087 56899
rect 25087 56865 25096 56899
rect 25044 56856 25096 56865
rect 25228 56856 25280 56908
rect 27068 56899 27120 56908
rect 22652 56788 22704 56840
rect 23756 56831 23808 56840
rect 23756 56797 23765 56831
rect 23765 56797 23799 56831
rect 23799 56797 23808 56831
rect 24216 56831 24268 56840
rect 23756 56788 23808 56797
rect 24216 56797 24226 56831
rect 24226 56797 24268 56831
rect 24216 56788 24268 56797
rect 25136 56831 25188 56840
rect 25136 56797 25145 56831
rect 25145 56797 25179 56831
rect 25179 56797 25188 56831
rect 25596 56831 25648 56840
rect 25136 56788 25188 56797
rect 25596 56797 25606 56831
rect 25606 56797 25648 56831
rect 25596 56788 25648 56797
rect 26332 56831 26384 56840
rect 26332 56797 26341 56831
rect 26341 56797 26375 56831
rect 26375 56797 26384 56831
rect 26332 56788 26384 56797
rect 26424 56831 26476 56840
rect 26424 56797 26433 56831
rect 26433 56797 26467 56831
rect 26467 56797 26476 56831
rect 27068 56865 27077 56899
rect 27077 56865 27111 56899
rect 27111 56865 27120 56899
rect 27068 56856 27120 56865
rect 27620 56856 27672 56908
rect 26424 56788 26476 56797
rect 27528 56831 27580 56840
rect 27528 56797 27540 56831
rect 27540 56797 27574 56831
rect 27574 56797 27580 56831
rect 27804 56856 27856 56908
rect 27528 56788 27580 56797
rect 27988 56788 28040 56840
rect 28540 56856 28592 56908
rect 33048 56856 33100 56908
rect 33692 56924 33744 56976
rect 36268 56924 36320 56976
rect 41144 56924 41196 56976
rect 28724 56831 28776 56840
rect 28724 56797 28733 56831
rect 28733 56797 28767 56831
rect 28767 56797 28776 56831
rect 28724 56788 28776 56797
rect 28816 56788 28868 56840
rect 7288 56720 7340 56772
rect 16948 56652 17000 56704
rect 24032 56652 24084 56704
rect 24768 56652 24820 56704
rect 25688 56652 25740 56704
rect 26148 56695 26200 56704
rect 26148 56661 26157 56695
rect 26157 56661 26191 56695
rect 26191 56661 26200 56695
rect 26148 56652 26200 56661
rect 28632 56720 28684 56772
rect 28908 56720 28960 56772
rect 29552 56831 29604 56840
rect 29552 56797 29561 56831
rect 29561 56797 29595 56831
rect 29595 56797 29604 56831
rect 29736 56831 29788 56840
rect 29552 56788 29604 56797
rect 29736 56797 29745 56831
rect 29745 56797 29779 56831
rect 29779 56797 29788 56831
rect 29736 56788 29788 56797
rect 31668 56788 31720 56840
rect 32312 56831 32364 56840
rect 32312 56797 32321 56831
rect 32321 56797 32355 56831
rect 32355 56797 32364 56831
rect 32312 56788 32364 56797
rect 33876 56856 33928 56908
rect 33692 56831 33744 56840
rect 33692 56797 33701 56831
rect 33701 56797 33735 56831
rect 33735 56797 33744 56831
rect 33692 56788 33744 56797
rect 33784 56831 33836 56840
rect 33784 56797 33793 56831
rect 33793 56797 33827 56831
rect 33827 56797 33836 56831
rect 35624 56856 35676 56908
rect 38384 56856 38436 56908
rect 38660 56856 38712 56908
rect 41236 56856 41288 56908
rect 43352 56924 43404 56976
rect 43720 56924 43772 56976
rect 50620 56924 50672 56976
rect 43904 56899 43956 56908
rect 33784 56788 33836 56797
rect 35992 56831 36044 56840
rect 35992 56797 36001 56831
rect 36001 56797 36035 56831
rect 36035 56797 36044 56831
rect 35992 56788 36044 56797
rect 36268 56831 36320 56840
rect 36268 56797 36277 56831
rect 36277 56797 36311 56831
rect 36311 56797 36320 56831
rect 36268 56788 36320 56797
rect 36636 56788 36688 56840
rect 36820 56831 36872 56840
rect 36820 56797 36829 56831
rect 36829 56797 36863 56831
rect 36863 56797 36872 56831
rect 36820 56788 36872 56797
rect 37556 56788 37608 56840
rect 38016 56831 38068 56840
rect 38016 56797 38025 56831
rect 38025 56797 38059 56831
rect 38059 56797 38068 56831
rect 38016 56788 38068 56797
rect 38108 56831 38160 56840
rect 38108 56797 38117 56831
rect 38117 56797 38151 56831
rect 38151 56797 38160 56831
rect 38108 56788 38160 56797
rect 38752 56788 38804 56840
rect 39028 56788 39080 56840
rect 39856 56788 39908 56840
rect 40776 56788 40828 56840
rect 40960 56788 41012 56840
rect 41512 56788 41564 56840
rect 41788 56831 41840 56840
rect 41788 56797 41797 56831
rect 41797 56797 41831 56831
rect 41831 56797 41840 56831
rect 41788 56788 41840 56797
rect 43904 56865 43913 56899
rect 43913 56865 43947 56899
rect 43947 56865 43956 56899
rect 43904 56856 43956 56865
rect 48320 56856 48372 56908
rect 41972 56788 42024 56840
rect 43168 56788 43220 56840
rect 43352 56831 43404 56840
rect 43352 56797 43361 56831
rect 43361 56797 43395 56831
rect 43395 56797 43404 56831
rect 43352 56788 43404 56797
rect 43628 56788 43680 56840
rect 44088 56831 44140 56840
rect 44088 56797 44097 56831
rect 44097 56797 44131 56831
rect 44131 56797 44140 56831
rect 44088 56788 44140 56797
rect 44456 56831 44508 56840
rect 44456 56797 44465 56831
rect 44465 56797 44499 56831
rect 44499 56797 44508 56831
rect 44456 56788 44508 56797
rect 45192 56831 45244 56840
rect 34428 56720 34480 56772
rect 35808 56720 35860 56772
rect 42248 56720 42300 56772
rect 45192 56797 45201 56831
rect 45201 56797 45235 56831
rect 45235 56797 45244 56831
rect 45192 56788 45244 56797
rect 45836 56831 45888 56840
rect 45836 56797 45845 56831
rect 45845 56797 45879 56831
rect 45879 56797 45888 56831
rect 45836 56788 45888 56797
rect 48688 56831 48740 56840
rect 48688 56797 48697 56831
rect 48697 56797 48731 56831
rect 48731 56797 48740 56831
rect 48688 56788 48740 56797
rect 45008 56720 45060 56772
rect 54116 56720 54168 56772
rect 26516 56652 26568 56704
rect 29552 56652 29604 56704
rect 30840 56652 30892 56704
rect 32036 56652 32088 56704
rect 33232 56695 33284 56704
rect 33232 56661 33241 56695
rect 33241 56661 33275 56695
rect 33275 56661 33284 56695
rect 33232 56652 33284 56661
rect 34520 56652 34572 56704
rect 39488 56652 39540 56704
rect 40960 56695 41012 56704
rect 40960 56661 40969 56695
rect 40969 56661 41003 56695
rect 41003 56661 41012 56695
rect 40960 56652 41012 56661
rect 41144 56695 41196 56704
rect 41144 56661 41153 56695
rect 41153 56661 41187 56695
rect 41187 56661 41196 56695
rect 41144 56652 41196 56661
rect 41972 56652 42024 56704
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 23756 56448 23808 56500
rect 22560 56312 22612 56364
rect 24216 56355 24268 56364
rect 24216 56321 24225 56355
rect 24225 56321 24259 56355
rect 24259 56321 24268 56355
rect 25596 56448 25648 56500
rect 26240 56380 26292 56432
rect 24216 56312 24268 56321
rect 24492 56244 24544 56296
rect 24860 56244 24912 56296
rect 25872 56312 25924 56364
rect 26424 56312 26476 56364
rect 27896 56380 27948 56432
rect 28264 56423 28316 56432
rect 28264 56389 28273 56423
rect 28273 56389 28307 56423
rect 28307 56389 28316 56423
rect 28264 56380 28316 56389
rect 28724 56448 28776 56500
rect 28908 56448 28960 56500
rect 32220 56448 32272 56500
rect 33784 56448 33836 56500
rect 35532 56491 35584 56500
rect 35532 56457 35541 56491
rect 35541 56457 35575 56491
rect 35575 56457 35584 56491
rect 35532 56448 35584 56457
rect 36820 56448 36872 56500
rect 39488 56448 39540 56500
rect 35348 56380 35400 56432
rect 28816 56312 28868 56364
rect 29000 56312 29052 56364
rect 31668 56312 31720 56364
rect 32220 56355 32272 56364
rect 32220 56321 32229 56355
rect 32229 56321 32263 56355
rect 32263 56321 32272 56355
rect 33232 56355 33284 56364
rect 32220 56312 32272 56321
rect 27344 56287 27396 56296
rect 27344 56253 27353 56287
rect 27353 56253 27387 56287
rect 27387 56253 27396 56287
rect 27344 56244 27396 56253
rect 27988 56244 28040 56296
rect 29828 56287 29880 56296
rect 29828 56253 29837 56287
rect 29837 56253 29871 56287
rect 29871 56253 29880 56287
rect 29828 56244 29880 56253
rect 30840 56244 30892 56296
rect 24584 56108 24636 56160
rect 26608 56108 26660 56160
rect 27528 56176 27580 56228
rect 28724 56176 28776 56228
rect 29368 56108 29420 56160
rect 29736 56176 29788 56228
rect 31116 56176 31168 56228
rect 32772 56244 32824 56296
rect 33232 56321 33241 56355
rect 33241 56321 33275 56355
rect 33275 56321 33284 56355
rect 33232 56312 33284 56321
rect 34152 56355 34204 56364
rect 34152 56321 34161 56355
rect 34161 56321 34195 56355
rect 34195 56321 34204 56355
rect 34152 56312 34204 56321
rect 34428 56355 34480 56364
rect 34428 56321 34437 56355
rect 34437 56321 34471 56355
rect 34471 56321 34480 56355
rect 37464 56380 37516 56432
rect 38200 56380 38252 56432
rect 38844 56380 38896 56432
rect 35624 56355 35676 56364
rect 34428 56312 34480 56321
rect 33324 56244 33376 56296
rect 31208 56108 31260 56160
rect 32496 56108 32548 56160
rect 33416 56151 33468 56160
rect 33416 56117 33425 56151
rect 33425 56117 33459 56151
rect 33459 56117 33468 56151
rect 33416 56108 33468 56117
rect 33876 56244 33928 56296
rect 34336 56287 34388 56296
rect 34336 56253 34345 56287
rect 34345 56253 34379 56287
rect 34379 56253 34388 56287
rect 35624 56321 35633 56355
rect 35633 56321 35667 56355
rect 35667 56321 35676 56355
rect 35624 56312 35676 56321
rect 35808 56355 35860 56364
rect 35808 56321 35817 56355
rect 35817 56321 35851 56355
rect 35851 56321 35860 56355
rect 35808 56312 35860 56321
rect 35992 56355 36044 56364
rect 35992 56321 36001 56355
rect 36001 56321 36035 56355
rect 36035 56321 36044 56355
rect 35992 56312 36044 56321
rect 36452 56312 36504 56364
rect 37924 56312 37976 56364
rect 40132 56448 40184 56500
rect 40500 56448 40552 56500
rect 41880 56448 41932 56500
rect 42892 56448 42944 56500
rect 44272 56491 44324 56500
rect 44272 56457 44281 56491
rect 44281 56457 44315 56491
rect 44315 56457 44324 56491
rect 44272 56448 44324 56457
rect 45008 56448 45060 56500
rect 49700 56448 49752 56500
rect 51448 56491 51500 56500
rect 51448 56457 51457 56491
rect 51457 56457 51491 56491
rect 51491 56457 51500 56491
rect 51448 56448 51500 56457
rect 52828 56491 52880 56500
rect 52828 56457 52837 56491
rect 52837 56457 52871 56491
rect 52871 56457 52880 56491
rect 52828 56448 52880 56457
rect 53840 56491 53892 56500
rect 53840 56457 53849 56491
rect 53849 56457 53883 56491
rect 53883 56457 53892 56491
rect 53840 56448 53892 56457
rect 43996 56380 44048 56432
rect 39948 56355 40000 56364
rect 39948 56321 39957 56355
rect 39957 56321 39991 56355
rect 39991 56321 40000 56355
rect 39948 56312 40000 56321
rect 40132 56312 40184 56364
rect 41144 56355 41196 56364
rect 41144 56321 41153 56355
rect 41153 56321 41187 56355
rect 41187 56321 41196 56355
rect 41144 56312 41196 56321
rect 41972 56312 42024 56364
rect 44088 56355 44140 56364
rect 34336 56244 34388 56253
rect 34704 56244 34756 56296
rect 35716 56244 35768 56296
rect 38200 56244 38252 56296
rect 38752 56244 38804 56296
rect 40224 56287 40276 56296
rect 40224 56253 40233 56287
rect 40233 56253 40267 56287
rect 40267 56253 40276 56287
rect 40224 56244 40276 56253
rect 41512 56244 41564 56296
rect 43352 56287 43404 56296
rect 33600 56176 33652 56228
rect 34704 56108 34756 56160
rect 37372 56176 37424 56228
rect 38108 56219 38160 56228
rect 38108 56185 38117 56219
rect 38117 56185 38151 56219
rect 38151 56185 38160 56219
rect 38108 56176 38160 56185
rect 41880 56219 41932 56228
rect 41880 56185 41889 56219
rect 41889 56185 41923 56219
rect 41923 56185 41932 56219
rect 41880 56176 41932 56185
rect 42064 56176 42116 56228
rect 40408 56108 40460 56160
rect 40960 56108 41012 56160
rect 42248 56151 42300 56160
rect 42248 56117 42257 56151
rect 42257 56117 42291 56151
rect 42291 56117 42300 56151
rect 42248 56108 42300 56117
rect 43352 56253 43361 56287
rect 43361 56253 43395 56287
rect 43395 56253 43404 56287
rect 43352 56244 43404 56253
rect 44088 56321 44097 56355
rect 44097 56321 44131 56355
rect 44131 56321 44140 56355
rect 44088 56312 44140 56321
rect 45008 56312 45060 56364
rect 45284 56355 45336 56364
rect 45284 56321 45293 56355
rect 45293 56321 45327 56355
rect 45327 56321 45336 56355
rect 45284 56312 45336 56321
rect 46480 56312 46532 56364
rect 47400 56312 47452 56364
rect 48780 56312 48832 56364
rect 49240 56312 49292 56364
rect 44272 56244 44324 56296
rect 44640 56244 44692 56296
rect 42800 56176 42852 56228
rect 43260 56176 43312 56228
rect 42708 56108 42760 56160
rect 44364 56108 44416 56160
rect 44548 56108 44600 56160
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 23940 55947 23992 55956
rect 23940 55913 23949 55947
rect 23949 55913 23983 55947
rect 23983 55913 23992 55947
rect 23940 55904 23992 55913
rect 25136 55904 25188 55956
rect 25780 55904 25832 55956
rect 28264 55904 28316 55956
rect 29000 55904 29052 55956
rect 35440 55904 35492 55956
rect 37188 55904 37240 55956
rect 37464 55904 37516 55956
rect 38016 55904 38068 55956
rect 38292 55904 38344 55956
rect 40960 55904 41012 55956
rect 44272 55947 44324 55956
rect 26700 55836 26752 55888
rect 27896 55836 27948 55888
rect 28724 55836 28776 55888
rect 24584 55743 24636 55752
rect 24584 55709 24593 55743
rect 24593 55709 24627 55743
rect 24627 55709 24636 55743
rect 24584 55700 24636 55709
rect 29276 55768 29328 55820
rect 31576 55836 31628 55888
rect 33048 55879 33100 55888
rect 33048 55845 33057 55879
rect 33057 55845 33091 55879
rect 33091 55845 33100 55879
rect 33048 55836 33100 55845
rect 31300 55768 31352 55820
rect 31668 55811 31720 55820
rect 31668 55777 31677 55811
rect 31677 55777 31711 55811
rect 31711 55777 31720 55811
rect 31668 55768 31720 55777
rect 28816 55743 28868 55752
rect 28816 55709 28825 55743
rect 28825 55709 28859 55743
rect 28859 55709 28868 55743
rect 28816 55700 28868 55709
rect 28908 55743 28960 55752
rect 28908 55709 28917 55743
rect 28917 55709 28951 55743
rect 28951 55709 28960 55743
rect 28908 55700 28960 55709
rect 29736 55700 29788 55752
rect 30288 55743 30340 55752
rect 30288 55709 30297 55743
rect 30297 55709 30331 55743
rect 30331 55709 30340 55743
rect 30288 55700 30340 55709
rect 31944 55700 31996 55752
rect 32404 55700 32456 55752
rect 32588 55743 32640 55752
rect 32588 55709 32597 55743
rect 32597 55709 32631 55743
rect 32631 55709 32640 55743
rect 32588 55700 32640 55709
rect 33692 55836 33744 55888
rect 34060 55836 34112 55888
rect 36544 55836 36596 55888
rect 36912 55836 36964 55888
rect 35532 55768 35584 55820
rect 36084 55768 36136 55820
rect 27988 55675 28040 55684
rect 24492 55564 24544 55616
rect 27988 55641 27997 55675
rect 27997 55641 28031 55675
rect 28031 55641 28040 55675
rect 27988 55632 28040 55641
rect 29000 55632 29052 55684
rect 30104 55675 30156 55684
rect 30104 55641 30113 55675
rect 30113 55641 30147 55675
rect 30147 55641 30156 55675
rect 30104 55632 30156 55641
rect 29276 55564 29328 55616
rect 31852 55632 31904 55684
rect 32496 55675 32548 55684
rect 32496 55641 32505 55675
rect 32505 55641 32539 55675
rect 32539 55641 32548 55675
rect 33784 55700 33836 55752
rect 34336 55743 34388 55752
rect 34336 55709 34344 55743
rect 34344 55709 34378 55743
rect 34378 55709 34388 55743
rect 34336 55700 34388 55709
rect 34704 55700 34756 55752
rect 36268 55700 36320 55752
rect 36820 55743 36872 55752
rect 36820 55709 36829 55743
rect 36829 55709 36863 55743
rect 36863 55709 36872 55743
rect 36820 55700 36872 55709
rect 39672 55768 39724 55820
rect 32496 55632 32548 55641
rect 32772 55564 32824 55616
rect 35716 55632 35768 55684
rect 38200 55700 38252 55752
rect 38752 55700 38804 55752
rect 34520 55564 34572 55616
rect 34796 55564 34848 55616
rect 36084 55564 36136 55616
rect 36728 55607 36780 55616
rect 36728 55573 36737 55607
rect 36737 55573 36771 55607
rect 36771 55573 36780 55607
rect 36728 55564 36780 55573
rect 38476 55632 38528 55684
rect 39212 55700 39264 55752
rect 41328 55836 41380 55888
rect 44272 55913 44281 55947
rect 44281 55913 44315 55947
rect 44315 55913 44324 55947
rect 44272 55904 44324 55913
rect 44732 55904 44784 55956
rect 45100 55904 45152 55956
rect 47584 55947 47636 55956
rect 47584 55913 47593 55947
rect 47593 55913 47627 55947
rect 47627 55913 47636 55947
rect 47584 55904 47636 55913
rect 48320 55947 48372 55956
rect 48320 55913 48329 55947
rect 48329 55913 48363 55947
rect 48363 55913 48372 55947
rect 48320 55904 48372 55913
rect 41052 55768 41104 55820
rect 43628 55879 43680 55888
rect 43628 55845 43637 55879
rect 43637 55845 43671 55879
rect 43671 55845 43680 55879
rect 43628 55836 43680 55845
rect 40868 55743 40920 55752
rect 40868 55709 40877 55743
rect 40877 55709 40911 55743
rect 40911 55709 40920 55743
rect 40868 55700 40920 55709
rect 40960 55700 41012 55752
rect 43260 55768 43312 55820
rect 39304 55675 39356 55684
rect 39304 55641 39313 55675
rect 39313 55641 39347 55675
rect 39347 55641 39356 55675
rect 39304 55632 39356 55641
rect 41972 55700 42024 55752
rect 43444 55743 43496 55752
rect 43444 55709 43453 55743
rect 43453 55709 43487 55743
rect 43487 55709 43496 55743
rect 44088 55768 44140 55820
rect 44364 55768 44416 55820
rect 45284 55768 45336 55820
rect 43444 55700 43496 55709
rect 43720 55743 43772 55752
rect 43720 55709 43729 55743
rect 43729 55709 43763 55743
rect 43763 55709 43772 55743
rect 44548 55743 44600 55752
rect 43720 55700 43772 55709
rect 44548 55709 44557 55743
rect 44557 55709 44591 55743
rect 44591 55709 44600 55743
rect 44548 55700 44600 55709
rect 43352 55632 43404 55684
rect 44456 55675 44508 55684
rect 44456 55641 44465 55675
rect 44465 55641 44499 55675
rect 44499 55641 44508 55675
rect 44456 55632 44508 55641
rect 39028 55564 39080 55616
rect 39764 55564 39816 55616
rect 40960 55564 41012 55616
rect 41512 55564 41564 55616
rect 46756 55564 46808 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 25044 55360 25096 55412
rect 25964 55403 26016 55412
rect 25964 55369 25973 55403
rect 25973 55369 26007 55403
rect 26007 55369 26016 55403
rect 25964 55360 26016 55369
rect 26976 55360 27028 55412
rect 27252 55360 27304 55412
rect 29092 55360 29144 55412
rect 29368 55292 29420 55344
rect 25504 55267 25556 55276
rect 25504 55233 25513 55267
rect 25513 55233 25547 55267
rect 25547 55233 25556 55267
rect 25504 55224 25556 55233
rect 26148 55267 26200 55276
rect 26148 55233 26157 55267
rect 26157 55233 26191 55267
rect 26191 55233 26200 55267
rect 26148 55224 26200 55233
rect 26608 55267 26660 55276
rect 26608 55233 26617 55267
rect 26617 55233 26651 55267
rect 26651 55233 26660 55267
rect 26608 55224 26660 55233
rect 26976 55224 27028 55276
rect 28816 55156 28868 55208
rect 29552 55267 29604 55276
rect 29552 55233 29561 55267
rect 29561 55233 29595 55267
rect 29595 55233 29604 55267
rect 31392 55292 31444 55344
rect 31576 55360 31628 55412
rect 35716 55360 35768 55412
rect 35808 55360 35860 55412
rect 37924 55403 37976 55412
rect 37924 55369 37933 55403
rect 37933 55369 37967 55403
rect 37967 55369 37976 55403
rect 37924 55360 37976 55369
rect 38476 55360 38528 55412
rect 40868 55360 40920 55412
rect 41788 55403 41840 55412
rect 41788 55369 41797 55403
rect 41797 55369 41831 55403
rect 41831 55369 41840 55403
rect 41788 55360 41840 55369
rect 31852 55292 31904 55344
rect 34244 55292 34296 55344
rect 29552 55224 29604 55233
rect 30012 55224 30064 55276
rect 30472 55224 30524 55276
rect 30932 55267 30984 55276
rect 30932 55233 30941 55267
rect 30941 55233 30975 55267
rect 30975 55233 30984 55267
rect 30932 55224 30984 55233
rect 31116 55267 31168 55276
rect 31116 55233 31125 55267
rect 31125 55233 31159 55267
rect 31159 55233 31168 55267
rect 31116 55224 31168 55233
rect 31760 55224 31812 55276
rect 32772 55224 32824 55276
rect 34520 55267 34572 55276
rect 34520 55233 34529 55267
rect 34529 55233 34563 55267
rect 34563 55233 34572 55267
rect 34520 55224 34572 55233
rect 35440 55335 35492 55344
rect 35440 55301 35449 55335
rect 35449 55301 35483 55335
rect 35483 55301 35492 55335
rect 35440 55292 35492 55301
rect 37556 55292 37608 55344
rect 37372 55267 37424 55276
rect 32404 55156 32456 55208
rect 34244 55156 34296 55208
rect 35992 55156 36044 55208
rect 37372 55233 37381 55267
rect 37381 55233 37415 55267
rect 37415 55233 37424 55267
rect 37372 55224 37424 55233
rect 38016 55224 38068 55276
rect 38752 55292 38804 55344
rect 38936 55292 38988 55344
rect 43168 55360 43220 55412
rect 45284 55360 45336 55412
rect 54208 55360 54260 55412
rect 39212 55224 39264 55276
rect 39580 55224 39632 55276
rect 40040 55224 40092 55276
rect 42064 55267 42116 55276
rect 42064 55233 42073 55267
rect 42073 55233 42107 55267
rect 42107 55233 42116 55267
rect 42064 55224 42116 55233
rect 37280 55156 37332 55208
rect 38752 55156 38804 55208
rect 28908 55088 28960 55140
rect 31300 55088 31352 55140
rect 32588 55088 32640 55140
rect 34428 55088 34480 55140
rect 34704 55131 34756 55140
rect 34704 55097 34713 55131
rect 34713 55097 34747 55131
rect 34747 55097 34756 55131
rect 41696 55156 41748 55208
rect 43720 55292 43772 55344
rect 43444 55224 43496 55276
rect 44180 55224 44232 55276
rect 42432 55199 42484 55208
rect 42432 55165 42441 55199
rect 42441 55165 42475 55199
rect 42475 55165 42484 55199
rect 42432 55156 42484 55165
rect 34704 55088 34756 55097
rect 39120 55088 39172 55140
rect 39304 55088 39356 55140
rect 43628 55088 43680 55140
rect 24584 55063 24636 55072
rect 24584 55029 24593 55063
rect 24593 55029 24627 55063
rect 24627 55029 24636 55063
rect 24584 55020 24636 55029
rect 32036 55063 32088 55072
rect 32036 55029 32045 55063
rect 32045 55029 32079 55063
rect 32079 55029 32088 55063
rect 32036 55020 32088 55029
rect 32404 55063 32456 55072
rect 32404 55029 32413 55063
rect 32413 55029 32447 55063
rect 32447 55029 32456 55063
rect 32404 55020 32456 55029
rect 33048 55063 33100 55072
rect 33048 55029 33057 55063
rect 33057 55029 33091 55063
rect 33091 55029 33100 55063
rect 33048 55020 33100 55029
rect 33600 55020 33652 55072
rect 33968 55020 34020 55072
rect 39580 55020 39632 55072
rect 40408 55020 40460 55072
rect 41052 55020 41104 55072
rect 41880 55020 41932 55072
rect 42064 55020 42116 55072
rect 43260 55020 43312 55072
rect 45928 55156 45980 55208
rect 44916 55063 44968 55072
rect 44916 55029 44925 55063
rect 44925 55029 44959 55063
rect 44959 55029 44968 55063
rect 44916 55020 44968 55029
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 25320 54816 25372 54868
rect 28080 54816 28132 54868
rect 28356 54859 28408 54868
rect 28356 54825 28365 54859
rect 28365 54825 28399 54859
rect 28399 54825 28408 54859
rect 28356 54816 28408 54825
rect 30472 54816 30524 54868
rect 31116 54816 31168 54868
rect 29276 54748 29328 54800
rect 29644 54748 29696 54800
rect 33324 54816 33376 54868
rect 36544 54859 36596 54868
rect 36544 54825 36553 54859
rect 36553 54825 36587 54859
rect 36587 54825 36596 54859
rect 36544 54816 36596 54825
rect 37188 54859 37240 54868
rect 37188 54825 37197 54859
rect 37197 54825 37231 54859
rect 37231 54825 37240 54859
rect 37188 54816 37240 54825
rect 38200 54816 38252 54868
rect 38936 54859 38988 54868
rect 38936 54825 38945 54859
rect 38945 54825 38979 54859
rect 38979 54825 38988 54859
rect 38936 54816 38988 54825
rect 40132 54859 40184 54868
rect 40132 54825 40141 54859
rect 40141 54825 40175 54859
rect 40175 54825 40184 54859
rect 40132 54816 40184 54825
rect 41972 54816 42024 54868
rect 42892 54859 42944 54868
rect 42892 54825 42901 54859
rect 42901 54825 42935 54859
rect 42935 54825 42944 54859
rect 42892 54816 42944 54825
rect 43536 54859 43588 54868
rect 43536 54825 43545 54859
rect 43545 54825 43579 54859
rect 43579 54825 43588 54859
rect 43536 54816 43588 54825
rect 31760 54748 31812 54800
rect 28632 54680 28684 54732
rect 29092 54723 29144 54732
rect 29092 54689 29101 54723
rect 29101 54689 29135 54723
rect 29135 54689 29144 54723
rect 29092 54680 29144 54689
rect 30104 54680 30156 54732
rect 28540 54612 28592 54664
rect 29368 54612 29420 54664
rect 32404 54723 32456 54732
rect 31300 54612 31352 54664
rect 32404 54689 32413 54723
rect 32413 54689 32447 54723
rect 32447 54689 32456 54723
rect 32404 54680 32456 54689
rect 33416 54748 33468 54800
rect 33048 54612 33100 54664
rect 34520 54680 34572 54732
rect 34612 54680 34664 54732
rect 34980 54680 35032 54732
rect 33968 54655 34020 54664
rect 33968 54621 33977 54655
rect 33977 54621 34011 54655
rect 34011 54621 34020 54655
rect 33968 54612 34020 54621
rect 34428 54612 34480 54664
rect 34704 54612 34756 54664
rect 33508 54544 33560 54596
rect 34888 54544 34940 54596
rect 35900 54612 35952 54664
rect 38568 54748 38620 54800
rect 42800 54748 42852 54800
rect 38384 54723 38436 54732
rect 38384 54689 38393 54723
rect 38393 54689 38427 54723
rect 38427 54689 38436 54723
rect 40868 54723 40920 54732
rect 38384 54680 38436 54689
rect 39120 54655 39172 54664
rect 39120 54621 39129 54655
rect 39129 54621 39163 54655
rect 39163 54621 39172 54655
rect 39120 54612 39172 54621
rect 39212 54655 39264 54664
rect 39212 54621 39221 54655
rect 39221 54621 39255 54655
rect 39255 54621 39264 54655
rect 39212 54612 39264 54621
rect 39580 54612 39632 54664
rect 38752 54544 38804 54596
rect 39764 54587 39816 54596
rect 39764 54553 39773 54587
rect 39773 54553 39807 54587
rect 39807 54553 39816 54587
rect 39764 54544 39816 54553
rect 40868 54689 40877 54723
rect 40877 54689 40911 54723
rect 40911 54689 40920 54723
rect 40868 54680 40920 54689
rect 40960 54655 41012 54664
rect 40960 54621 40969 54655
rect 40969 54621 41003 54655
rect 41003 54621 41012 54655
rect 40960 54612 41012 54621
rect 41788 54655 41840 54664
rect 41788 54621 41797 54655
rect 41797 54621 41831 54655
rect 41831 54621 41840 54655
rect 41788 54612 41840 54621
rect 41880 54655 41932 54664
rect 41880 54621 41889 54655
rect 41889 54621 41923 54655
rect 41923 54621 41932 54655
rect 41880 54612 41932 54621
rect 43168 54612 43220 54664
rect 44916 54544 44968 54596
rect 24584 54519 24636 54528
rect 24584 54485 24593 54519
rect 24593 54485 24627 54519
rect 24627 54485 24636 54519
rect 26424 54519 26476 54528
rect 24584 54476 24636 54485
rect 26424 54485 26433 54519
rect 26433 54485 26467 54519
rect 26467 54485 26476 54519
rect 26424 54476 26476 54485
rect 30012 54476 30064 54528
rect 30472 54476 30524 54528
rect 33140 54476 33192 54528
rect 34428 54476 34480 54528
rect 42248 54476 42300 54528
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 25872 54315 25924 54324
rect 25872 54281 25881 54315
rect 25881 54281 25915 54315
rect 25915 54281 25924 54315
rect 25872 54272 25924 54281
rect 27620 54272 27672 54324
rect 29552 54315 29604 54324
rect 29552 54281 29561 54315
rect 29561 54281 29595 54315
rect 29595 54281 29604 54315
rect 29552 54272 29604 54281
rect 31116 54272 31168 54324
rect 32772 54272 32824 54324
rect 33508 54315 33560 54324
rect 33508 54281 33517 54315
rect 33517 54281 33551 54315
rect 33551 54281 33560 54315
rect 33508 54272 33560 54281
rect 33692 54272 33744 54324
rect 37372 54272 37424 54324
rect 39580 54315 39632 54324
rect 39580 54281 39589 54315
rect 39589 54281 39623 54315
rect 39623 54281 39632 54315
rect 39580 54272 39632 54281
rect 40408 54272 40460 54324
rect 41880 54272 41932 54324
rect 42064 54272 42116 54324
rect 42708 54272 42760 54324
rect 30012 54204 30064 54256
rect 30472 54247 30524 54256
rect 30472 54213 30481 54247
rect 30481 54213 30515 54247
rect 30515 54213 30524 54247
rect 30472 54204 30524 54213
rect 31944 54204 31996 54256
rect 29000 54136 29052 54188
rect 30104 54136 30156 54188
rect 30932 54179 30984 54188
rect 30932 54145 30941 54179
rect 30941 54145 30975 54179
rect 30975 54145 30984 54179
rect 30932 54136 30984 54145
rect 33600 54204 33652 54256
rect 37464 54204 37516 54256
rect 38384 54247 38436 54256
rect 38384 54213 38393 54247
rect 38393 54213 38427 54247
rect 38427 54213 38436 54247
rect 38384 54204 38436 54213
rect 38568 54247 38620 54256
rect 38568 54213 38577 54247
rect 38577 54213 38611 54247
rect 38611 54213 38620 54247
rect 38568 54204 38620 54213
rect 39948 54204 40000 54256
rect 32404 54136 32456 54188
rect 34244 54136 34296 54188
rect 34704 54179 34756 54188
rect 34704 54145 34713 54179
rect 34713 54145 34747 54179
rect 34747 54145 34756 54179
rect 34704 54136 34756 54145
rect 34980 54179 35032 54188
rect 34980 54145 34989 54179
rect 34989 54145 35023 54179
rect 35023 54145 35032 54179
rect 34980 54136 35032 54145
rect 35624 54179 35676 54188
rect 35624 54145 35633 54179
rect 35633 54145 35667 54179
rect 35667 54145 35676 54179
rect 35624 54136 35676 54145
rect 36084 54179 36136 54188
rect 36084 54145 36093 54179
rect 36093 54145 36127 54179
rect 36127 54145 36136 54179
rect 36084 54136 36136 54145
rect 36360 54136 36412 54188
rect 39672 54136 39724 54188
rect 40316 54136 40368 54188
rect 40776 54136 40828 54188
rect 41696 54136 41748 54188
rect 42432 54136 42484 54188
rect 34888 54111 34940 54120
rect 34888 54077 34897 54111
rect 34897 54077 34931 54111
rect 34931 54077 34940 54111
rect 34888 54068 34940 54077
rect 26424 54000 26476 54052
rect 27344 54000 27396 54052
rect 28172 54000 28224 54052
rect 29368 54043 29420 54052
rect 29368 54009 29377 54043
rect 29377 54009 29411 54043
rect 29411 54009 29420 54043
rect 29368 54000 29420 54009
rect 31668 54000 31720 54052
rect 40224 54068 40276 54120
rect 32036 53932 32088 53984
rect 40040 53932 40092 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 28172 53771 28224 53780
rect 28172 53737 28181 53771
rect 28181 53737 28215 53771
rect 28215 53737 28224 53771
rect 28172 53728 28224 53737
rect 29184 53728 29236 53780
rect 29920 53728 29972 53780
rect 32772 53728 32824 53780
rect 33600 53771 33652 53780
rect 33600 53737 33609 53771
rect 33609 53737 33643 53771
rect 33643 53737 33652 53771
rect 33600 53728 33652 53737
rect 34428 53728 34480 53780
rect 35624 53728 35676 53780
rect 35900 53728 35952 53780
rect 37740 53728 37792 53780
rect 38844 53728 38896 53780
rect 39856 53728 39908 53780
rect 39948 53728 40000 53780
rect 40776 53771 40828 53780
rect 37464 53660 37516 53712
rect 40776 53737 40785 53771
rect 40785 53737 40819 53771
rect 40819 53737 40828 53771
rect 40776 53728 40828 53737
rect 42708 53728 42760 53780
rect 29276 53567 29328 53576
rect 29276 53533 29285 53567
rect 29285 53533 29319 53567
rect 29319 53533 29328 53567
rect 29276 53524 29328 53533
rect 29368 53524 29420 53576
rect 30288 53524 30340 53576
rect 31392 53524 31444 53576
rect 31944 53431 31996 53440
rect 31944 53397 31953 53431
rect 31953 53397 31987 53431
rect 31987 53397 31996 53431
rect 31944 53388 31996 53397
rect 33140 53567 33192 53576
rect 33140 53533 33149 53567
rect 33149 53533 33183 53567
rect 33183 53533 33192 53567
rect 33140 53524 33192 53533
rect 36084 53524 36136 53576
rect 39948 53524 40000 53576
rect 34152 53456 34204 53508
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 30288 53227 30340 53236
rect 30288 53193 30297 53227
rect 30297 53193 30331 53227
rect 30331 53193 30340 53227
rect 30288 53184 30340 53193
rect 31944 53184 31996 53236
rect 35624 53184 35676 53236
rect 38660 53184 38712 53236
rect 39948 53227 40000 53236
rect 39948 53193 39957 53227
rect 39957 53193 39991 53227
rect 39991 53193 40000 53227
rect 39948 53184 40000 53193
rect 33784 53116 33836 53168
rect 36452 53116 36504 53168
rect 29460 53048 29512 53100
rect 36084 53091 36136 53100
rect 36084 53057 36093 53091
rect 36093 53057 36127 53091
rect 36127 53057 36136 53091
rect 36084 53048 36136 53057
rect 34520 53023 34572 53032
rect 34520 52989 34529 53023
rect 34529 52989 34563 53023
rect 34563 52989 34572 53023
rect 34520 52980 34572 52989
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 29368 52683 29420 52692
rect 29368 52649 29377 52683
rect 29377 52649 29411 52683
rect 29411 52649 29420 52683
rect 29368 52640 29420 52649
rect 35624 52640 35676 52692
rect 36176 52640 36228 52692
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 26424 8075 26476 8084
rect 26424 8041 26433 8075
rect 26433 8041 26467 8075
rect 26467 8041 26476 8075
rect 26424 8032 26476 8041
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 24952 7420 25004 7472
rect 30288 7352 30340 7404
rect 22560 7284 22612 7336
rect 26792 7327 26844 7336
rect 26792 7293 26801 7327
rect 26801 7293 26835 7327
rect 26835 7293 26844 7327
rect 26792 7284 26844 7293
rect 26700 7148 26752 7200
rect 29736 7191 29788 7200
rect 29736 7157 29745 7191
rect 29745 7157 29779 7191
rect 29779 7157 29788 7191
rect 29736 7148 29788 7157
rect 30380 7191 30432 7200
rect 30380 7157 30389 7191
rect 30389 7157 30423 7191
rect 30423 7157 30432 7191
rect 30380 7148 30432 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 25596 6808 25648 6860
rect 28632 6851 28684 6860
rect 28632 6817 28641 6851
rect 28641 6817 28675 6851
rect 28675 6817 28684 6851
rect 28632 6808 28684 6817
rect 26608 6740 26660 6792
rect 29552 6740 29604 6792
rect 31024 6783 31076 6792
rect 31024 6749 31033 6783
rect 31033 6749 31067 6783
rect 31067 6749 31076 6783
rect 31024 6740 31076 6749
rect 31760 6740 31812 6792
rect 26516 6715 26568 6724
rect 26516 6681 26525 6715
rect 26525 6681 26559 6715
rect 26559 6681 26568 6715
rect 28172 6715 28224 6724
rect 26516 6672 26568 6681
rect 24860 6604 24912 6656
rect 26884 6604 26936 6656
rect 28172 6681 28181 6715
rect 28181 6681 28215 6715
rect 28215 6681 28224 6715
rect 28172 6672 28224 6681
rect 30380 6604 30432 6656
rect 32220 6647 32272 6656
rect 32220 6613 32229 6647
rect 32229 6613 32263 6647
rect 32263 6613 32272 6647
rect 32220 6604 32272 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 29736 6375 29788 6384
rect 29736 6341 29745 6375
rect 29745 6341 29779 6375
rect 29779 6341 29788 6375
rect 29736 6332 29788 6341
rect 38200 6332 38252 6384
rect 24492 6264 24544 6316
rect 26608 6264 26660 6316
rect 29552 6307 29604 6316
rect 29552 6273 29561 6307
rect 29561 6273 29595 6307
rect 29595 6273 29604 6307
rect 29552 6264 29604 6273
rect 26240 6196 26292 6248
rect 27896 6239 27948 6248
rect 27896 6205 27905 6239
rect 27905 6205 27939 6239
rect 27939 6205 27948 6239
rect 27896 6196 27948 6205
rect 30196 6239 30248 6248
rect 30196 6205 30205 6239
rect 30205 6205 30239 6239
rect 30239 6205 30248 6239
rect 30196 6196 30248 6205
rect 30288 6196 30340 6248
rect 34428 6239 34480 6248
rect 34428 6205 34437 6239
rect 34437 6205 34471 6239
rect 34471 6205 34480 6239
rect 34428 6196 34480 6205
rect 37924 6196 37976 6248
rect 23940 6060 23992 6112
rect 24676 6060 24728 6112
rect 31208 6060 31260 6112
rect 33048 6103 33100 6112
rect 33048 6069 33057 6103
rect 33057 6069 33091 6103
rect 33091 6069 33100 6103
rect 33048 6060 33100 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 24676 5763 24728 5772
rect 24676 5729 24685 5763
rect 24685 5729 24719 5763
rect 24719 5729 24728 5763
rect 24676 5720 24728 5729
rect 24860 5763 24912 5772
rect 24860 5729 24869 5763
rect 24869 5729 24903 5763
rect 24903 5729 24912 5763
rect 24860 5720 24912 5729
rect 26148 5763 26200 5772
rect 26148 5729 26157 5763
rect 26157 5729 26191 5763
rect 26191 5729 26200 5763
rect 26148 5720 26200 5729
rect 28080 5763 28132 5772
rect 28080 5729 28089 5763
rect 28089 5729 28123 5763
rect 28123 5729 28132 5763
rect 28080 5720 28132 5729
rect 30104 5720 30156 5772
rect 30288 5763 30340 5772
rect 30288 5729 30297 5763
rect 30297 5729 30331 5763
rect 30331 5729 30340 5763
rect 30288 5720 30340 5729
rect 31024 5763 31076 5772
rect 31024 5729 31033 5763
rect 31033 5729 31067 5763
rect 31067 5729 31076 5763
rect 31024 5720 31076 5729
rect 31208 5763 31260 5772
rect 31208 5729 31217 5763
rect 31217 5729 31251 5763
rect 31251 5729 31260 5763
rect 31208 5720 31260 5729
rect 31668 5763 31720 5772
rect 31668 5729 31677 5763
rect 31677 5729 31711 5763
rect 31711 5729 31720 5763
rect 31668 5720 31720 5729
rect 23112 5652 23164 5704
rect 24492 5652 24544 5704
rect 26056 5652 26108 5704
rect 26516 5652 26568 5704
rect 27528 5695 27580 5704
rect 27528 5661 27537 5695
rect 27537 5661 27571 5695
rect 27571 5661 27580 5695
rect 27528 5652 27580 5661
rect 30380 5652 30432 5704
rect 33140 5652 33192 5704
rect 26976 5584 27028 5636
rect 31024 5584 31076 5636
rect 31760 5584 31812 5636
rect 35348 5652 35400 5704
rect 24124 5559 24176 5568
rect 24124 5525 24133 5559
rect 24133 5525 24167 5559
rect 24167 5525 24176 5559
rect 24124 5516 24176 5525
rect 33232 5516 33284 5568
rect 34796 5516 34848 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 26976 5312 27028 5364
rect 24124 5244 24176 5296
rect 26884 5287 26936 5296
rect 26884 5253 26893 5287
rect 26893 5253 26927 5287
rect 26927 5253 26936 5287
rect 26884 5244 26936 5253
rect 34796 5287 34848 5296
rect 34796 5253 34805 5287
rect 34805 5253 34839 5287
rect 34839 5253 34848 5287
rect 34796 5244 34848 5253
rect 24492 5176 24544 5228
rect 22284 5108 22336 5160
rect 25412 5108 25464 5160
rect 26056 5176 26108 5228
rect 26700 5219 26752 5228
rect 26700 5185 26709 5219
rect 26709 5185 26743 5219
rect 26743 5185 26752 5219
rect 26700 5176 26752 5185
rect 28356 5151 28408 5160
rect 28356 5117 28365 5151
rect 28365 5117 28399 5151
rect 28399 5117 28408 5151
rect 28356 5108 28408 5117
rect 30288 5151 30340 5160
rect 30288 5117 30297 5151
rect 30297 5117 30331 5151
rect 30331 5117 30340 5151
rect 30288 5108 30340 5117
rect 30564 5151 30616 5160
rect 30564 5117 30573 5151
rect 30573 5117 30607 5151
rect 30607 5117 30616 5151
rect 30564 5108 30616 5117
rect 33324 5151 33376 5160
rect 33324 5117 33333 5151
rect 33333 5117 33367 5151
rect 33367 5117 33376 5151
rect 33324 5108 33376 5117
rect 22836 4972 22888 5024
rect 31024 4972 31076 5024
rect 35900 4972 35952 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 22560 4811 22612 4820
rect 22560 4777 22569 4811
rect 22569 4777 22603 4811
rect 22603 4777 22612 4811
rect 22560 4768 22612 4777
rect 27528 4811 27580 4820
rect 27528 4777 27537 4811
rect 27537 4777 27571 4811
rect 27571 4777 27580 4811
rect 27528 4768 27580 4777
rect 23388 4700 23440 4752
rect 19340 4607 19392 4616
rect 19340 4573 19349 4607
rect 19349 4573 19383 4607
rect 19383 4573 19392 4607
rect 19340 4564 19392 4573
rect 20352 4564 20404 4616
rect 21732 4564 21784 4616
rect 22192 4564 22244 4616
rect 24492 4632 24544 4684
rect 30012 4675 30064 4684
rect 30012 4641 30021 4675
rect 30021 4641 30055 4675
rect 30055 4641 30064 4675
rect 30012 4632 30064 4641
rect 31760 4632 31812 4684
rect 33140 4700 33192 4752
rect 37280 4700 37332 4752
rect 32220 4675 32272 4684
rect 32220 4641 32229 4675
rect 32229 4641 32263 4675
rect 32263 4641 32272 4675
rect 32220 4632 32272 4641
rect 32772 4675 32824 4684
rect 32772 4641 32781 4675
rect 32781 4641 32815 4675
rect 32815 4641 32824 4675
rect 32772 4632 32824 4641
rect 31024 4607 31076 4616
rect 31024 4573 31033 4607
rect 31033 4573 31067 4607
rect 31067 4573 31076 4607
rect 31024 4564 31076 4573
rect 36820 4607 36872 4616
rect 36820 4573 36829 4607
rect 36829 4573 36863 4607
rect 36863 4573 36872 4607
rect 36820 4564 36872 4573
rect 37464 4564 37516 4616
rect 38936 4607 38988 4616
rect 38936 4573 38945 4607
rect 38945 4573 38979 4607
rect 38979 4573 38988 4607
rect 38936 4564 38988 4573
rect 27528 4496 27580 4548
rect 29460 4496 29512 4548
rect 34980 4539 35032 4548
rect 34980 4505 34989 4539
rect 34989 4505 35023 4539
rect 35023 4505 35032 4539
rect 34980 4496 35032 4505
rect 37372 4496 37424 4548
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 30288 4224 30340 4276
rect 22284 4131 22336 4140
rect 22284 4097 22293 4131
rect 22293 4097 22327 4131
rect 22327 4097 22336 4131
rect 22284 4088 22336 4097
rect 25596 4131 25648 4140
rect 25596 4097 25605 4131
rect 25605 4097 25639 4131
rect 25639 4097 25648 4131
rect 25596 4088 25648 4097
rect 26240 4131 26292 4140
rect 26240 4097 26249 4131
rect 26249 4097 26283 4131
rect 26283 4097 26292 4131
rect 26240 4088 26292 4097
rect 29552 4088 29604 4140
rect 30104 4088 30156 4140
rect 33048 4131 33100 4140
rect 33048 4097 33057 4131
rect 33057 4097 33091 4131
rect 33091 4097 33100 4131
rect 33048 4088 33100 4097
rect 35348 4131 35400 4140
rect 35348 4097 35357 4131
rect 35357 4097 35391 4131
rect 35391 4097 35400 4131
rect 35348 4088 35400 4097
rect 36820 4088 36872 4140
rect 20628 4020 20680 4072
rect 22744 4063 22796 4072
rect 22744 4029 22753 4063
rect 22753 4029 22787 4063
rect 22787 4029 22796 4063
rect 22744 4020 22796 4029
rect 22928 4063 22980 4072
rect 22928 4029 22937 4063
rect 22937 4029 22971 4063
rect 22971 4029 22980 4063
rect 22928 4020 22980 4029
rect 16304 3884 16356 3936
rect 17592 3884 17644 3936
rect 18420 3884 18472 3936
rect 19432 3884 19484 3936
rect 22008 3952 22060 4004
rect 24492 3884 24544 3936
rect 27436 4020 27488 4072
rect 29736 4020 29788 4072
rect 30656 4063 30708 4072
rect 30656 4029 30665 4063
rect 30665 4029 30699 4063
rect 30699 4029 30708 4063
rect 30656 4020 30708 4029
rect 31392 4063 31444 4072
rect 27988 3952 28040 4004
rect 31392 4029 31401 4063
rect 31401 4029 31435 4063
rect 31435 4029 31444 4063
rect 31392 4020 31444 4029
rect 33232 4063 33284 4072
rect 33232 4029 33241 4063
rect 33241 4029 33275 4063
rect 33275 4029 33284 4063
rect 33232 4020 33284 4029
rect 37004 4063 37056 4072
rect 33048 3952 33100 4004
rect 37004 4029 37013 4063
rect 37013 4029 37047 4063
rect 37047 4029 37056 4063
rect 37004 4020 37056 4029
rect 37188 4063 37240 4072
rect 37188 4029 37197 4063
rect 37197 4029 37231 4063
rect 37231 4029 37240 4063
rect 37188 4020 37240 4029
rect 34152 3952 34204 4004
rect 27252 3884 27304 3936
rect 33876 3884 33928 3936
rect 34980 3884 35032 3936
rect 35440 3927 35492 3936
rect 35440 3893 35449 3927
rect 35449 3893 35483 3927
rect 35483 3893 35492 3927
rect 35440 3884 35492 3893
rect 39120 3952 39172 4004
rect 37740 3884 37792 3936
rect 40224 3884 40276 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 22744 3680 22796 3732
rect 27436 3723 27488 3732
rect 27436 3689 27445 3723
rect 27445 3689 27479 3723
rect 27479 3689 27488 3723
rect 27436 3680 27488 3689
rect 27988 3723 28040 3732
rect 27988 3689 27997 3723
rect 27997 3689 28031 3723
rect 28031 3689 28040 3723
rect 27988 3680 28040 3689
rect 30656 3680 30708 3732
rect 37372 3723 37424 3732
rect 37372 3689 37381 3723
rect 37381 3689 37415 3723
rect 37415 3689 37424 3723
rect 37372 3680 37424 3689
rect 37924 3723 37976 3732
rect 37924 3689 37933 3723
rect 37933 3689 37967 3723
rect 37967 3689 37976 3723
rect 37924 3680 37976 3689
rect 38108 3680 38160 3732
rect 21456 3612 21508 3664
rect 20076 3544 20128 3596
rect 26976 3612 27028 3664
rect 29184 3612 29236 3664
rect 32220 3612 32272 3664
rect 29644 3544 29696 3596
rect 32496 3587 32548 3596
rect 32496 3553 32505 3587
rect 32505 3553 32539 3587
rect 32539 3553 32548 3587
rect 32496 3544 32548 3553
rect 35348 3544 35400 3596
rect 36636 3612 36688 3664
rect 39396 3612 39448 3664
rect 42156 3612 42208 3664
rect 43260 3612 43312 3664
rect 45468 3612 45520 3664
rect 35532 3544 35584 3596
rect 9312 3476 9364 3528
rect 10232 3476 10284 3528
rect 11888 3476 11940 3528
rect 12716 3476 12768 3528
rect 13544 3476 13596 3528
rect 14372 3476 14424 3528
rect 14924 3476 14976 3528
rect 15752 3476 15804 3528
rect 16856 3476 16908 3528
rect 17868 3476 17920 3528
rect 18144 3476 18196 3528
rect 22560 3519 22612 3528
rect 22560 3485 22569 3519
rect 22569 3485 22603 3519
rect 22603 3485 22612 3519
rect 22560 3476 22612 3485
rect 24584 3476 24636 3528
rect 26516 3519 26568 3528
rect 26516 3485 26525 3519
rect 26525 3485 26559 3519
rect 26559 3485 26568 3519
rect 26516 3476 26568 3485
rect 27436 3476 27488 3528
rect 33692 3519 33744 3528
rect 33692 3485 33701 3519
rect 33701 3485 33735 3519
rect 33735 3485 33744 3519
rect 34336 3519 34388 3528
rect 33692 3476 33744 3485
rect 34336 3485 34345 3519
rect 34345 3485 34379 3519
rect 34379 3485 34388 3519
rect 34336 3476 34388 3485
rect 34980 3519 35032 3528
rect 34980 3485 34989 3519
rect 34989 3485 35023 3519
rect 35023 3485 35032 3519
rect 34980 3476 35032 3485
rect 37372 3476 37424 3528
rect 38568 3544 38620 3596
rect 40776 3544 40828 3596
rect 44088 3544 44140 3596
rect 23848 3408 23900 3460
rect 26332 3451 26384 3460
rect 26332 3417 26341 3451
rect 26341 3417 26375 3451
rect 26375 3417 26384 3451
rect 26332 3408 26384 3417
rect 29092 3408 29144 3460
rect 31024 3408 31076 3460
rect 35348 3408 35400 3460
rect 36912 3408 36964 3460
rect 39028 3408 39080 3460
rect 23664 3340 23716 3392
rect 34796 3340 34848 3392
rect 38752 3340 38804 3392
rect 41328 3476 41380 3528
rect 42708 3476 42760 3528
rect 44916 3476 44968 3528
rect 46296 3476 46348 3528
rect 47124 3476 47176 3528
rect 47676 3476 47728 3528
rect 49056 3476 49108 3528
rect 49608 3476 49660 3528
rect 50988 3476 51040 3528
rect 51540 3476 51592 3528
rect 40040 3340 40092 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 24952 3136 25004 3188
rect 29460 3179 29512 3188
rect 29460 3145 29469 3179
rect 29469 3145 29503 3179
rect 29503 3145 29512 3179
rect 29460 3136 29512 3145
rect 36360 3136 36412 3188
rect 37464 3136 37516 3188
rect 19984 3068 20036 3120
rect 24216 3068 24268 3120
rect 35440 3068 35492 3120
rect 37556 3068 37608 3120
rect 38108 3068 38160 3120
rect 21180 3000 21232 3052
rect 22192 3000 22244 3052
rect 22560 3000 22612 3052
rect 24584 3043 24636 3052
rect 24584 3009 24593 3043
rect 24593 3009 24627 3043
rect 24627 3009 24636 3043
rect 24584 3000 24636 3009
rect 26516 3000 26568 3052
rect 29552 3043 29604 3052
rect 29552 3009 29561 3043
rect 29561 3009 29595 3043
rect 29595 3009 29604 3043
rect 29552 3000 29604 3009
rect 34980 3000 35032 3052
rect 16028 2932 16080 2984
rect 18972 2932 19024 2984
rect 19524 2864 19576 2916
rect 19984 2907 20036 2916
rect 19984 2873 19993 2907
rect 19993 2873 20027 2907
rect 20027 2873 20036 2907
rect 19984 2864 20036 2873
rect 7656 2796 7708 2848
rect 8208 2796 8260 2848
rect 8944 2796 8996 2848
rect 9956 2796 10008 2848
rect 10508 2796 10560 2848
rect 11060 2796 11112 2848
rect 11612 2796 11664 2848
rect 12164 2796 12216 2848
rect 12992 2796 13044 2848
rect 13820 2796 13872 2848
rect 14096 2839 14148 2848
rect 14096 2805 14105 2839
rect 14105 2805 14139 2839
rect 14139 2805 14148 2839
rect 14096 2796 14148 2805
rect 15200 2796 15252 2848
rect 16580 2796 16632 2848
rect 17316 2796 17368 2848
rect 22560 2864 22612 2916
rect 25228 2932 25280 2984
rect 27804 2932 27856 2984
rect 29460 2932 29512 2984
rect 28908 2864 28960 2916
rect 31116 2932 31168 2984
rect 30380 2864 30432 2916
rect 30840 2864 30892 2916
rect 31944 2932 31996 2984
rect 34704 2975 34756 2984
rect 34704 2941 34713 2975
rect 34713 2941 34747 2975
rect 34747 2941 34756 2975
rect 34704 2932 34756 2941
rect 34520 2864 34572 2916
rect 25044 2796 25096 2848
rect 25412 2796 25464 2848
rect 26424 2796 26476 2848
rect 33600 2796 33652 2848
rect 35808 2864 35860 2916
rect 38384 3000 38436 3052
rect 41052 3000 41104 3052
rect 39672 2932 39724 2984
rect 41880 2932 41932 2984
rect 44364 2932 44416 2984
rect 46572 2932 46624 2984
rect 49884 2932 49936 2984
rect 52092 2932 52144 2984
rect 35440 2796 35492 2848
rect 35900 2796 35952 2848
rect 38016 2864 38068 2916
rect 38936 2864 38988 2916
rect 39028 2864 39080 2916
rect 40500 2864 40552 2916
rect 42984 2864 43036 2916
rect 45192 2864 45244 2916
rect 47400 2864 47452 2916
rect 48780 2864 48832 2916
rect 50712 2864 50764 2916
rect 43628 2796 43680 2848
rect 45744 2796 45796 2848
rect 47952 2796 48004 2848
rect 49332 2796 49384 2848
rect 51264 2796 51316 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 22928 2592 22980 2644
rect 23848 2592 23900 2644
rect 25228 2635 25280 2644
rect 25228 2601 25237 2635
rect 25237 2601 25271 2635
rect 25271 2601 25280 2635
rect 25228 2592 25280 2601
rect 26332 2592 26384 2644
rect 27804 2635 27856 2644
rect 27804 2601 27813 2635
rect 27813 2601 27847 2635
rect 27847 2601 27856 2635
rect 27804 2592 27856 2601
rect 29092 2635 29144 2644
rect 29092 2601 29101 2635
rect 29101 2601 29135 2635
rect 29135 2601 29144 2635
rect 29092 2592 29144 2601
rect 29644 2635 29696 2644
rect 29644 2601 29653 2635
rect 29653 2601 29687 2635
rect 29687 2601 29696 2635
rect 29644 2592 29696 2601
rect 30380 2635 30432 2644
rect 30380 2601 30389 2635
rect 30389 2601 30423 2635
rect 30423 2601 30432 2635
rect 30380 2592 30432 2601
rect 31116 2635 31168 2644
rect 31116 2601 31125 2635
rect 31125 2601 31159 2635
rect 31159 2601 31168 2635
rect 31116 2592 31168 2601
rect 33692 2592 33744 2644
rect 34704 2592 34756 2644
rect 35348 2592 35400 2644
rect 37004 2592 37056 2644
rect 38200 2635 38252 2644
rect 38200 2601 38209 2635
rect 38209 2601 38243 2635
rect 38243 2601 38252 2635
rect 38200 2592 38252 2601
rect 38752 2635 38804 2644
rect 38752 2601 38761 2635
rect 38761 2601 38795 2635
rect 38795 2601 38804 2635
rect 38752 2592 38804 2601
rect 40040 2635 40092 2644
rect 40040 2601 40049 2635
rect 40049 2601 40083 2635
rect 40083 2601 40092 2635
rect 40040 2592 40092 2601
rect 8576 2524 8628 2576
rect 12440 2524 12492 2576
rect 18696 2524 18748 2576
rect 25596 2524 25648 2576
rect 34520 2524 34572 2576
rect 37188 2524 37240 2576
rect 39948 2524 40000 2576
rect 43812 2524 43864 2576
rect 46848 2524 46900 2576
rect 51816 2524 51868 2576
rect 10784 2456 10836 2508
rect 14648 2456 14700 2508
rect 17132 2456 17184 2508
rect 20904 2456 20956 2508
rect 25872 2456 25924 2508
rect 38844 2456 38896 2508
rect 42432 2456 42484 2508
rect 44640 2456 44692 2508
rect 48228 2456 48280 2508
rect 50160 2456 50212 2508
rect 52368 2456 52420 2508
rect 9680 2388 9732 2440
rect 11336 2388 11388 2440
rect 13268 2388 13320 2440
rect 15476 2388 15528 2440
rect 19984 2388 20036 2440
rect 23296 2388 23348 2440
rect 22284 2320 22336 2372
rect 27436 2388 27488 2440
rect 29552 2388 29604 2440
rect 34336 2388 34388 2440
rect 37372 2388 37424 2440
rect 19340 2252 19392 2304
rect 19524 2252 19576 2304
rect 22192 2252 22244 2304
rect 28172 2320 28224 2372
rect 36084 2320 36136 2372
rect 41604 2320 41656 2372
rect 46020 2388 46072 2440
rect 48504 2388 48556 2440
rect 50620 2388 50672 2440
rect 23296 2252 23348 2304
rect 25320 2252 25372 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 19984 2048 20036 2100
rect 24768 2048 24820 2100
<< metal2 >>
rect 3698 59200 3754 60000
rect 4158 59200 4214 60000
rect 4618 59200 4674 60000
rect 5078 59200 5134 60000
rect 5538 59200 5594 60000
rect 5998 59200 6054 60000
rect 6458 59200 6514 60000
rect 6918 59200 6974 60000
rect 7378 59200 7434 60000
rect 7838 59200 7894 60000
rect 8298 59200 8354 60000
rect 8758 59200 8814 60000
rect 9218 59200 9274 60000
rect 9678 59200 9734 60000
rect 10138 59200 10194 60000
rect 10598 59200 10654 60000
rect 10704 59214 11008 59242
rect 3712 57526 3740 59200
rect 3700 57520 3752 57526
rect 3700 57462 3752 57468
rect 3712 57050 3740 57462
rect 4632 57458 4660 59200
rect 5092 57594 5120 59200
rect 5080 57588 5132 57594
rect 5080 57530 5132 57536
rect 4620 57452 4672 57458
rect 4620 57394 4672 57400
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 6012 57050 6040 59200
rect 6472 57458 6500 59200
rect 6460 57452 6512 57458
rect 6460 57394 6512 57400
rect 7288 57384 7340 57390
rect 7288 57326 7340 57332
rect 7300 57254 7328 57326
rect 7288 57248 7340 57254
rect 7288 57190 7340 57196
rect 3700 57044 3752 57050
rect 3700 56986 3752 56992
rect 6000 57044 6052 57050
rect 6000 56986 6052 56992
rect 7300 56778 7328 57190
rect 7392 57050 7420 59200
rect 7852 57458 7880 59200
rect 8772 57458 8800 59200
rect 9232 57458 9260 59200
rect 10152 57458 10180 59200
rect 10612 59106 10640 59200
rect 10704 59106 10732 59214
rect 10612 59078 10732 59106
rect 10980 57610 11008 59214
rect 11058 59200 11114 60000
rect 11518 59200 11574 60000
rect 11978 59200 12034 60000
rect 12438 59200 12494 60000
rect 12898 59200 12954 60000
rect 13358 59200 13414 60000
rect 13818 59200 13874 60000
rect 14278 59200 14334 60000
rect 14738 59200 14794 60000
rect 15198 59200 15254 60000
rect 15658 59200 15714 60000
rect 16118 59200 16174 60000
rect 16578 59200 16634 60000
rect 17038 59200 17094 60000
rect 17498 59200 17554 60000
rect 17958 59200 18014 60000
rect 18418 59200 18474 60000
rect 18878 59200 18934 60000
rect 19338 59200 19394 60000
rect 19798 59200 19854 60000
rect 20258 59200 20314 60000
rect 20718 59200 20774 60000
rect 21178 59200 21234 60000
rect 21638 59200 21694 60000
rect 22098 59200 22154 60000
rect 22558 59200 22614 60000
rect 23018 59200 23074 60000
rect 23478 59200 23534 60000
rect 23938 59200 23994 60000
rect 24398 59200 24454 60000
rect 24858 59200 24914 60000
rect 25318 59200 25374 60000
rect 25778 59200 25834 60000
rect 26238 59200 26294 60000
rect 26698 59200 26754 60000
rect 27158 59200 27214 60000
rect 27618 59200 27674 60000
rect 28078 59200 28134 60000
rect 28538 59200 28594 60000
rect 28998 59200 29054 60000
rect 29458 59200 29514 60000
rect 29918 59200 29974 60000
rect 30378 59200 30434 60000
rect 30838 59200 30894 60000
rect 31298 59200 31354 60000
rect 31758 59200 31814 60000
rect 32218 59200 32274 60000
rect 32678 59200 32734 60000
rect 33138 59200 33194 60000
rect 33598 59200 33654 60000
rect 34058 59200 34114 60000
rect 34518 59200 34574 60000
rect 34978 59200 35034 60000
rect 35438 59200 35494 60000
rect 35898 59200 35954 60000
rect 36358 59200 36414 60000
rect 36818 59200 36874 60000
rect 37278 59200 37334 60000
rect 37738 59200 37794 60000
rect 38198 59200 38254 60000
rect 38658 59200 38714 60000
rect 39118 59200 39174 60000
rect 39578 59200 39634 60000
rect 40038 59200 40094 60000
rect 40144 59214 40356 59242
rect 10980 57594 11100 57610
rect 10980 57588 11112 57594
rect 10980 57582 11060 57588
rect 11060 57530 11112 57536
rect 7840 57452 7892 57458
rect 7840 57394 7892 57400
rect 8760 57452 8812 57458
rect 8760 57394 8812 57400
rect 9220 57452 9272 57458
rect 9220 57394 9272 57400
rect 10140 57452 10192 57458
rect 10140 57394 10192 57400
rect 11336 57452 11388 57458
rect 11336 57394 11388 57400
rect 7380 57044 7432 57050
rect 7380 56986 7432 56992
rect 11348 56914 11376 57394
rect 11532 57050 11560 59200
rect 11992 57594 12020 59200
rect 11980 57588 12032 57594
rect 11980 57530 12032 57536
rect 12346 57488 12402 57497
rect 12346 57423 12348 57432
rect 12400 57423 12402 57432
rect 12348 57394 12400 57400
rect 12912 57050 12940 59200
rect 13372 57594 13400 59200
rect 13360 57588 13412 57594
rect 13360 57530 13412 57536
rect 14292 57458 14320 59200
rect 14752 57594 14780 59200
rect 15200 57928 15252 57934
rect 15200 57870 15252 57876
rect 14740 57588 14792 57594
rect 14740 57530 14792 57536
rect 15212 57458 15240 57870
rect 15672 57458 15700 59200
rect 16132 57594 16160 59200
rect 16120 57588 16172 57594
rect 16120 57530 16172 57536
rect 14280 57452 14332 57458
rect 14280 57394 14332 57400
rect 15200 57452 15252 57458
rect 15200 57394 15252 57400
rect 15660 57452 15712 57458
rect 15660 57394 15712 57400
rect 16948 57316 17000 57322
rect 16948 57258 17000 57264
rect 11520 57044 11572 57050
rect 11520 56986 11572 56992
rect 12900 57044 12952 57050
rect 12900 56986 12952 56992
rect 11336 56908 11388 56914
rect 11336 56850 11388 56856
rect 7288 56772 7340 56778
rect 7288 56714 7340 56720
rect 16960 56710 16988 57258
rect 17052 57050 17080 59200
rect 17512 57594 17540 59200
rect 17500 57588 17552 57594
rect 17500 57530 17552 57536
rect 18432 57050 18460 59200
rect 18892 57594 18920 59200
rect 19812 58290 19840 59200
rect 19812 58262 20024 58290
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 18880 57588 18932 57594
rect 18880 57530 18932 57536
rect 19996 57458 20024 58262
rect 20272 57594 20300 59200
rect 20996 57792 21048 57798
rect 20996 57734 21048 57740
rect 20260 57588 20312 57594
rect 20260 57530 20312 57536
rect 21008 57458 21036 57734
rect 19248 57452 19300 57458
rect 19248 57394 19300 57400
rect 19984 57452 20036 57458
rect 19984 57394 20036 57400
rect 20996 57452 21048 57458
rect 20996 57394 21048 57400
rect 17040 57044 17092 57050
rect 17040 56986 17092 56992
rect 18420 57044 18472 57050
rect 18420 56986 18472 56992
rect 19260 56982 19288 57394
rect 21192 57050 21220 59200
rect 21652 57594 21680 59200
rect 22008 57860 22060 57866
rect 22008 57802 22060 57808
rect 21640 57588 21692 57594
rect 21640 57530 21692 57536
rect 22020 57458 22048 57802
rect 22008 57452 22060 57458
rect 22008 57394 22060 57400
rect 21364 57316 21416 57322
rect 21364 57258 21416 57264
rect 21180 57044 21232 57050
rect 21180 56986 21232 56992
rect 19248 56976 19300 56982
rect 19248 56918 19300 56924
rect 21376 56914 21404 57258
rect 22468 57248 22520 57254
rect 22468 57190 22520 57196
rect 22480 56982 22508 57190
rect 22468 56976 22520 56982
rect 22468 56918 22520 56924
rect 21364 56908 21416 56914
rect 21364 56850 21416 56856
rect 16948 56704 17000 56710
rect 16948 56646 17000 56652
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 22572 56370 22600 59200
rect 23032 57594 23060 59200
rect 23020 57588 23072 57594
rect 23020 57530 23072 57536
rect 23204 57520 23256 57526
rect 23204 57462 23256 57468
rect 22652 57248 22704 57254
rect 22652 57190 22704 57196
rect 22664 56846 22692 57190
rect 23216 57050 23244 57462
rect 23756 57452 23808 57458
rect 23756 57394 23808 57400
rect 23204 57044 23256 57050
rect 23204 56986 23256 56992
rect 23768 56846 23796 57394
rect 22652 56840 22704 56846
rect 22652 56782 22704 56788
rect 23756 56840 23808 56846
rect 23756 56782 23808 56788
rect 23768 56506 23796 56782
rect 23756 56500 23808 56506
rect 23756 56442 23808 56448
rect 22560 56364 22612 56370
rect 22560 56306 22612 56312
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 23952 55962 23980 59200
rect 24412 57594 24440 59200
rect 24676 57860 24728 57866
rect 24676 57802 24728 57808
rect 24768 57860 24820 57866
rect 24768 57802 24820 57808
rect 24688 57594 24716 57802
rect 24400 57588 24452 57594
rect 24400 57530 24452 57536
rect 24676 57588 24728 57594
rect 24676 57530 24728 57536
rect 24780 57458 24808 57802
rect 25044 57792 25096 57798
rect 25044 57734 25096 57740
rect 24768 57452 24820 57458
rect 24768 57394 24820 57400
rect 24032 56908 24084 56914
rect 24032 56850 24084 56856
rect 24044 56710 24072 56850
rect 24216 56840 24268 56846
rect 24216 56782 24268 56788
rect 24032 56704 24084 56710
rect 24032 56646 24084 56652
rect 24228 56370 24256 56782
rect 24780 56710 24808 57394
rect 25056 56914 25084 57734
rect 25228 57248 25280 57254
rect 25228 57190 25280 57196
rect 25240 56914 25268 57190
rect 24860 56908 24912 56914
rect 24860 56850 24912 56856
rect 25044 56908 25096 56914
rect 25044 56850 25096 56856
rect 25228 56908 25280 56914
rect 25228 56850 25280 56856
rect 24768 56704 24820 56710
rect 24768 56646 24820 56652
rect 24216 56364 24268 56370
rect 24216 56306 24268 56312
rect 24872 56302 24900 56850
rect 24492 56296 24544 56302
rect 24492 56238 24544 56244
rect 24860 56296 24912 56302
rect 24860 56238 24912 56244
rect 23940 55956 23992 55962
rect 23940 55898 23992 55904
rect 24504 55622 24532 56238
rect 24584 56160 24636 56166
rect 24584 56102 24636 56108
rect 24596 55758 24624 56102
rect 24584 55752 24636 55758
rect 24584 55694 24636 55700
rect 24492 55616 24544 55622
rect 24544 55564 24624 55570
rect 24492 55558 24624 55564
rect 24504 55542 24624 55558
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 24504 55493 24532 55542
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 24596 55078 24624 55542
rect 25056 55418 25084 56850
rect 25136 56840 25188 56846
rect 25136 56782 25188 56788
rect 25148 55962 25176 56782
rect 25136 55956 25188 55962
rect 25136 55898 25188 55904
rect 25044 55412 25096 55418
rect 25044 55354 25096 55360
rect 24584 55072 24636 55078
rect 24584 55014 24636 55020
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 24596 54534 24624 55014
rect 25332 54874 25360 59200
rect 25688 57928 25740 57934
rect 25688 57870 25740 57876
rect 25596 57452 25648 57458
rect 25596 57394 25648 57400
rect 25504 57248 25556 57254
rect 25504 57190 25556 57196
rect 25516 55282 25544 57190
rect 25608 56930 25636 57394
rect 25700 57050 25728 57870
rect 25688 57044 25740 57050
rect 25688 56986 25740 56992
rect 25608 56902 25728 56930
rect 25596 56840 25648 56846
rect 25596 56782 25648 56788
rect 25608 56506 25636 56782
rect 25700 56710 25728 56902
rect 25688 56704 25740 56710
rect 25688 56646 25740 56652
rect 25596 56500 25648 56506
rect 25596 56442 25648 56448
rect 25700 56273 25728 56646
rect 25686 56264 25742 56273
rect 25686 56199 25742 56208
rect 25792 55962 25820 59200
rect 25964 57588 26016 57594
rect 25964 57530 26016 57536
rect 25872 56364 25924 56370
rect 25872 56306 25924 56312
rect 25780 55956 25832 55962
rect 25780 55898 25832 55904
rect 25504 55276 25556 55282
rect 25504 55218 25556 55224
rect 25320 54868 25372 54874
rect 25320 54810 25372 54816
rect 24584 54528 24636 54534
rect 24584 54470 24636 54476
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 25884 54330 25912 56306
rect 25976 55418 26004 57530
rect 26424 57452 26476 57458
rect 26424 57394 26476 57400
rect 26148 57384 26200 57390
rect 26148 57326 26200 57332
rect 26160 56794 26188 57326
rect 26436 56846 26464 57394
rect 26332 56840 26384 56846
rect 26330 56808 26332 56817
rect 26424 56840 26476 56846
rect 26384 56808 26386 56817
rect 26160 56766 26280 56794
rect 26148 56704 26200 56710
rect 26148 56646 26200 56652
rect 25964 55412 26016 55418
rect 25964 55354 26016 55360
rect 26160 55282 26188 56646
rect 26252 56438 26280 56766
rect 26424 56782 26476 56788
rect 26514 56808 26570 56817
rect 26330 56743 26386 56752
rect 26240 56432 26292 56438
rect 26240 56374 26292 56380
rect 26436 56370 26464 56782
rect 26514 56743 26570 56752
rect 26528 56710 26556 56743
rect 26516 56704 26568 56710
rect 26516 56646 26568 56652
rect 26424 56364 26476 56370
rect 26424 56306 26476 56312
rect 26608 56160 26660 56166
rect 26608 56102 26660 56108
rect 26620 55282 26648 56102
rect 26712 55894 26740 59200
rect 27068 57588 27120 57594
rect 27068 57530 27120 57536
rect 26976 57044 27028 57050
rect 26976 56986 27028 56992
rect 26700 55888 26752 55894
rect 26700 55830 26752 55836
rect 26988 55418 27016 56986
rect 27080 56914 27108 57530
rect 27172 56930 27200 59200
rect 27620 57928 27672 57934
rect 27620 57870 27672 57876
rect 27632 57458 27660 57870
rect 27988 57792 28040 57798
rect 27988 57734 28040 57740
rect 27710 57488 27766 57497
rect 27620 57452 27672 57458
rect 27710 57423 27766 57432
rect 27896 57452 27948 57458
rect 27620 57394 27672 57400
rect 27724 57254 27752 57423
rect 27896 57394 27948 57400
rect 27712 57248 27764 57254
rect 27764 57208 27844 57236
rect 27712 57190 27764 57196
rect 27068 56908 27120 56914
rect 27172 56902 27292 56930
rect 27816 56914 27844 57208
rect 27068 56850 27120 56856
rect 27264 55418 27292 56902
rect 27620 56908 27672 56914
rect 27620 56850 27672 56856
rect 27804 56908 27856 56914
rect 27804 56850 27856 56856
rect 27528 56840 27580 56846
rect 27528 56782 27580 56788
rect 27344 56296 27396 56302
rect 27344 56238 27396 56244
rect 26976 55412 27028 55418
rect 26976 55354 27028 55360
rect 27252 55412 27304 55418
rect 27252 55354 27304 55360
rect 26988 55282 27016 55354
rect 26148 55276 26200 55282
rect 26148 55218 26200 55224
rect 26608 55276 26660 55282
rect 26608 55218 26660 55224
rect 26976 55276 27028 55282
rect 26976 55218 27028 55224
rect 26424 54528 26476 54534
rect 26424 54470 26476 54476
rect 25872 54324 25924 54330
rect 25872 54266 25924 54272
rect 26436 54058 26464 54470
rect 27356 54058 27384 56238
rect 27540 56234 27568 56782
rect 27528 56228 27580 56234
rect 27528 56170 27580 56176
rect 27632 54330 27660 56850
rect 27908 56438 27936 57394
rect 28000 56846 28028 57734
rect 27988 56840 28040 56846
rect 27988 56782 28040 56788
rect 27896 56432 27948 56438
rect 27896 56374 27948 56380
rect 27908 55894 27936 56374
rect 27988 56296 28040 56302
rect 27988 56238 28040 56244
rect 27896 55888 27948 55894
rect 27896 55830 27948 55836
rect 28000 55690 28028 56238
rect 27988 55684 28040 55690
rect 27988 55626 28040 55632
rect 28092 54874 28120 59200
rect 28552 57390 28580 59200
rect 28540 57384 28592 57390
rect 28540 57326 28592 57332
rect 28264 57316 28316 57322
rect 28264 57258 28316 57264
rect 28276 56438 28304 57258
rect 28356 57248 28408 57254
rect 28356 57190 28408 57196
rect 28264 56432 28316 56438
rect 28264 56374 28316 56380
rect 28276 55962 28304 56374
rect 28264 55956 28316 55962
rect 28264 55898 28316 55904
rect 28368 54874 28396 57190
rect 28540 56908 28592 56914
rect 28540 56850 28592 56856
rect 28080 54868 28132 54874
rect 28080 54810 28132 54816
rect 28356 54868 28408 54874
rect 28356 54810 28408 54816
rect 28552 54670 28580 56850
rect 28724 56840 28776 56846
rect 28724 56782 28776 56788
rect 28816 56840 28868 56846
rect 28816 56782 28868 56788
rect 28632 56772 28684 56778
rect 28632 56714 28684 56720
rect 28644 54738 28672 56714
rect 28736 56506 28764 56782
rect 28724 56500 28776 56506
rect 28724 56442 28776 56448
rect 28828 56370 28856 56782
rect 28908 56772 28960 56778
rect 28908 56714 28960 56720
rect 28920 56506 28948 56714
rect 29012 56522 29040 59200
rect 29184 57452 29236 57458
rect 29184 57394 29236 57400
rect 29276 57452 29328 57458
rect 29276 57394 29328 57400
rect 28908 56500 28960 56506
rect 29012 56494 29132 56522
rect 28908 56442 28960 56448
rect 28816 56364 28868 56370
rect 28816 56306 28868 56312
rect 29000 56364 29052 56370
rect 29000 56306 29052 56312
rect 28724 56228 28776 56234
rect 28724 56170 28776 56176
rect 28736 55894 28764 56170
rect 29012 55962 29040 56306
rect 29000 55956 29052 55962
rect 29000 55898 29052 55904
rect 28724 55888 28776 55894
rect 28724 55830 28776 55836
rect 28816 55752 28868 55758
rect 28816 55694 28868 55700
rect 28908 55752 28960 55758
rect 28908 55694 28960 55700
rect 28828 55214 28856 55694
rect 28816 55208 28868 55214
rect 28816 55150 28868 55156
rect 28920 55146 28948 55694
rect 29012 55690 29040 55898
rect 29000 55684 29052 55690
rect 29000 55626 29052 55632
rect 29104 55570 29132 56494
rect 29012 55542 29132 55570
rect 28908 55140 28960 55146
rect 28908 55082 28960 55088
rect 28632 54732 28684 54738
rect 28632 54674 28684 54680
rect 28540 54664 28592 54670
rect 28540 54606 28592 54612
rect 27620 54324 27672 54330
rect 27620 54266 27672 54272
rect 29012 54194 29040 55542
rect 29092 55412 29144 55418
rect 29092 55354 29144 55360
rect 29104 54738 29132 55354
rect 29092 54732 29144 54738
rect 29092 54674 29144 54680
rect 29000 54188 29052 54194
rect 29000 54130 29052 54136
rect 26424 54052 26476 54058
rect 26424 53994 26476 54000
rect 27344 54052 27396 54058
rect 27344 53994 27396 54000
rect 28172 54052 28224 54058
rect 28172 53994 28224 54000
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 26436 8090 26464 53994
rect 28184 53786 28212 53994
rect 29196 53786 29224 57394
rect 29288 56409 29316 57394
rect 29274 56400 29330 56409
rect 29274 56335 29330 56344
rect 29368 56160 29420 56166
rect 29368 56102 29420 56108
rect 29276 55820 29328 55826
rect 29276 55762 29328 55768
rect 29288 55622 29316 55762
rect 29276 55616 29328 55622
rect 29276 55558 29328 55564
rect 29380 55350 29408 56102
rect 29368 55344 29420 55350
rect 29368 55286 29420 55292
rect 29276 54800 29328 54806
rect 29276 54742 29328 54748
rect 28172 53780 28224 53786
rect 28172 53722 28224 53728
rect 29184 53780 29236 53786
rect 29184 53722 29236 53728
rect 29288 53582 29316 54742
rect 29368 54664 29420 54670
rect 29368 54606 29420 54612
rect 29380 54058 29408 54606
rect 29368 54052 29420 54058
rect 29368 53994 29420 54000
rect 29276 53576 29328 53582
rect 29276 53518 29328 53524
rect 29368 53576 29420 53582
rect 29368 53518 29420 53524
rect 29380 52698 29408 53518
rect 29472 53106 29500 59200
rect 29826 57080 29882 57089
rect 29826 57015 29828 57024
rect 29880 57015 29882 57024
rect 29828 56986 29880 56992
rect 29552 56840 29604 56846
rect 29736 56840 29788 56846
rect 29604 56800 29684 56828
rect 29552 56782 29604 56788
rect 29552 56704 29604 56710
rect 29550 56672 29552 56681
rect 29604 56672 29606 56681
rect 29550 56607 29606 56616
rect 29552 55276 29604 55282
rect 29552 55218 29604 55224
rect 29564 54330 29592 55218
rect 29656 54806 29684 56800
rect 29736 56782 29788 56788
rect 29748 56234 29776 56782
rect 29828 56296 29880 56302
rect 29828 56238 29880 56244
rect 29736 56228 29788 56234
rect 29736 56170 29788 56176
rect 29748 55758 29776 56170
rect 29840 56137 29868 56238
rect 29826 56128 29882 56137
rect 29826 56063 29882 56072
rect 29736 55752 29788 55758
rect 29736 55694 29788 55700
rect 29644 54800 29696 54806
rect 29644 54742 29696 54748
rect 29552 54324 29604 54330
rect 29552 54266 29604 54272
rect 29932 53786 29960 59200
rect 30012 57384 30064 57390
rect 30012 57326 30064 57332
rect 30024 57050 30052 57326
rect 30012 57044 30064 57050
rect 30012 56986 30064 56992
rect 30288 56976 30340 56982
rect 30288 56918 30340 56924
rect 30300 55758 30328 56918
rect 30392 56794 30420 59200
rect 30852 57050 30880 59200
rect 31312 57594 31340 59200
rect 31300 57588 31352 57594
rect 31300 57530 31352 57536
rect 31772 57458 31800 59200
rect 31392 57452 31444 57458
rect 31392 57394 31444 57400
rect 31760 57452 31812 57458
rect 31760 57394 31812 57400
rect 31208 57248 31260 57254
rect 31208 57190 31260 57196
rect 30840 57044 30892 57050
rect 30840 56986 30892 56992
rect 30392 56766 30512 56794
rect 30288 55752 30340 55758
rect 30288 55694 30340 55700
rect 30104 55684 30156 55690
rect 30104 55626 30156 55632
rect 30012 55276 30064 55282
rect 30012 55218 30064 55224
rect 30024 54534 30052 55218
rect 30116 54738 30144 55626
rect 30484 55282 30512 56766
rect 30840 56704 30892 56710
rect 30840 56646 30892 56652
rect 30852 56302 30880 56646
rect 30840 56296 30892 56302
rect 30840 56238 30892 56244
rect 31116 56228 31168 56234
rect 31116 56170 31168 56176
rect 31128 55808 31156 56170
rect 31220 56166 31248 57190
rect 31404 57050 31432 57394
rect 31668 57384 31720 57390
rect 31668 57326 31720 57332
rect 31392 57044 31444 57050
rect 31392 56986 31444 56992
rect 31680 56846 31708 57326
rect 32036 57248 32088 57254
rect 32036 57190 32088 57196
rect 31668 56840 31720 56846
rect 31668 56782 31720 56788
rect 31680 56370 31708 56782
rect 32048 56710 32076 57190
rect 32036 56704 32088 56710
rect 32036 56646 32088 56652
rect 31668 56364 31720 56370
rect 31668 56306 31720 56312
rect 31208 56160 31260 56166
rect 31208 56102 31260 56108
rect 31680 55944 31708 56306
rect 31680 55916 31800 55944
rect 31576 55888 31628 55894
rect 31576 55830 31628 55836
rect 31300 55820 31352 55826
rect 31128 55780 31300 55808
rect 31300 55762 31352 55768
rect 31588 55418 31616 55830
rect 31668 55820 31720 55826
rect 31668 55762 31720 55768
rect 31576 55412 31628 55418
rect 31576 55354 31628 55360
rect 31392 55344 31444 55350
rect 31392 55286 31444 55292
rect 30472 55276 30524 55282
rect 30472 55218 30524 55224
rect 30932 55276 30984 55282
rect 30932 55218 30984 55224
rect 31116 55276 31168 55282
rect 31116 55218 31168 55224
rect 30484 54874 30512 55218
rect 30472 54868 30524 54874
rect 30472 54810 30524 54816
rect 30104 54732 30156 54738
rect 30104 54674 30156 54680
rect 30012 54528 30064 54534
rect 30012 54470 30064 54476
rect 30024 54262 30052 54470
rect 30012 54256 30064 54262
rect 30012 54198 30064 54204
rect 30116 54194 30144 54674
rect 30472 54528 30524 54534
rect 30472 54470 30524 54476
rect 30484 54262 30512 54470
rect 30472 54256 30524 54262
rect 30472 54198 30524 54204
rect 30944 54194 30972 55218
rect 31128 54874 31156 55218
rect 31300 55140 31352 55146
rect 31300 55082 31352 55088
rect 31116 54868 31168 54874
rect 31116 54810 31168 54816
rect 31128 54330 31156 54810
rect 31312 54670 31340 55082
rect 31300 54664 31352 54670
rect 31300 54606 31352 54612
rect 31116 54324 31168 54330
rect 31116 54266 31168 54272
rect 30104 54188 30156 54194
rect 30104 54130 30156 54136
rect 30932 54188 30984 54194
rect 30932 54130 30984 54136
rect 29920 53780 29972 53786
rect 29920 53722 29972 53728
rect 31404 53582 31432 55286
rect 31680 54058 31708 55762
rect 31772 55282 31800 55916
rect 31944 55752 31996 55758
rect 31944 55694 31996 55700
rect 31852 55684 31904 55690
rect 31852 55626 31904 55632
rect 31864 55350 31892 55626
rect 31852 55344 31904 55350
rect 31852 55286 31904 55292
rect 31760 55276 31812 55282
rect 31760 55218 31812 55224
rect 31772 54806 31800 55218
rect 31760 54800 31812 54806
rect 31760 54742 31812 54748
rect 31956 54262 31984 55694
rect 32048 55078 32076 56646
rect 32232 56506 32260 59200
rect 32588 57384 32640 57390
rect 32588 57326 32640 57332
rect 32312 56840 32364 56846
rect 32310 56808 32312 56817
rect 32364 56808 32366 56817
rect 32310 56743 32366 56752
rect 32220 56500 32272 56506
rect 32220 56442 32272 56448
rect 32220 56364 32272 56370
rect 32220 56306 32272 56312
rect 32232 56137 32260 56306
rect 32496 56160 32548 56166
rect 32218 56128 32274 56137
rect 32496 56102 32548 56108
rect 32218 56063 32274 56072
rect 32404 55752 32456 55758
rect 32404 55694 32456 55700
rect 32416 55214 32444 55694
rect 32508 55690 32536 56102
rect 32600 55758 32628 57326
rect 32588 55752 32640 55758
rect 32588 55694 32640 55700
rect 32496 55684 32548 55690
rect 32496 55626 32548 55632
rect 32404 55208 32456 55214
rect 32404 55150 32456 55156
rect 32600 55146 32628 55694
rect 32692 55321 32720 59200
rect 33152 57390 33180 59200
rect 33140 57384 33192 57390
rect 33140 57326 33192 57332
rect 33048 56908 33100 56914
rect 33048 56850 33100 56856
rect 32772 56296 32824 56302
rect 32772 56238 32824 56244
rect 32784 55622 32812 56238
rect 33060 55894 33088 56850
rect 33232 56704 33284 56710
rect 33232 56646 33284 56652
rect 33244 56370 33272 56646
rect 33232 56364 33284 56370
rect 33232 56306 33284 56312
rect 33324 56296 33376 56302
rect 33324 56238 33376 56244
rect 33048 55888 33100 55894
rect 33048 55830 33100 55836
rect 32772 55616 32824 55622
rect 32772 55558 32824 55564
rect 32678 55312 32734 55321
rect 32678 55247 32734 55256
rect 32772 55276 32824 55282
rect 32772 55218 32824 55224
rect 32588 55140 32640 55146
rect 32588 55082 32640 55088
rect 32036 55072 32088 55078
rect 32036 55014 32088 55020
rect 32404 55072 32456 55078
rect 32404 55014 32456 55020
rect 31944 54256 31996 54262
rect 31944 54198 31996 54204
rect 31668 54052 31720 54058
rect 31668 53994 31720 54000
rect 30288 53576 30340 53582
rect 30288 53518 30340 53524
rect 31392 53576 31444 53582
rect 31392 53518 31444 53524
rect 30300 53242 30328 53518
rect 31956 53446 31984 54198
rect 32048 53990 32076 55014
rect 32416 54738 32444 55014
rect 32404 54732 32456 54738
rect 32404 54674 32456 54680
rect 32416 54194 32444 54674
rect 32784 54330 32812 55218
rect 33048 55072 33100 55078
rect 33048 55014 33100 55020
rect 33060 54670 33088 55014
rect 33336 54874 33364 56238
rect 33612 56234 33640 59200
rect 33692 57520 33744 57526
rect 33692 57462 33744 57468
rect 33704 56982 33732 57462
rect 33876 57248 33928 57254
rect 33876 57190 33928 57196
rect 33692 56976 33744 56982
rect 33692 56918 33744 56924
rect 33888 56914 33916 57190
rect 33876 56908 33928 56914
rect 33876 56850 33928 56856
rect 33692 56840 33744 56846
rect 33690 56808 33692 56817
rect 33784 56840 33836 56846
rect 33744 56808 33746 56817
rect 33784 56782 33836 56788
rect 33690 56743 33746 56752
rect 33600 56228 33652 56234
rect 33600 56170 33652 56176
rect 33416 56160 33468 56166
rect 33416 56102 33468 56108
rect 33324 54868 33376 54874
rect 33324 54810 33376 54816
rect 33428 54806 33456 56102
rect 33704 55894 33732 56743
rect 33796 56506 33824 56782
rect 33784 56500 33836 56506
rect 33784 56442 33836 56448
rect 33888 56302 33916 56850
rect 33876 56296 33928 56302
rect 33876 56238 33928 56244
rect 34072 55894 34100 59200
rect 34244 57588 34296 57594
rect 34244 57530 34296 57536
rect 34256 57050 34284 57530
rect 34532 57526 34560 59200
rect 34520 57520 34572 57526
rect 34520 57462 34572 57468
rect 34428 57316 34480 57322
rect 34428 57258 34480 57264
rect 34244 57044 34296 57050
rect 34244 56986 34296 56992
rect 34440 56778 34468 57258
rect 34612 57248 34664 57254
rect 34992 57236 35020 59200
rect 34612 57190 34664 57196
rect 34808 57208 35020 57236
rect 35348 57248 35400 57254
rect 34428 56772 34480 56778
rect 34428 56714 34480 56720
rect 34440 56370 34468 56714
rect 34520 56704 34572 56710
rect 34518 56672 34520 56681
rect 34572 56672 34574 56681
rect 34518 56607 34574 56616
rect 34152 56364 34204 56370
rect 34152 56306 34204 56312
rect 34428 56364 34480 56370
rect 34428 56306 34480 56312
rect 33692 55888 33744 55894
rect 33692 55830 33744 55836
rect 34060 55888 34112 55894
rect 34060 55830 34112 55836
rect 33600 55072 33652 55078
rect 33600 55014 33652 55020
rect 33416 54800 33468 54806
rect 33416 54742 33468 54748
rect 33048 54664 33100 54670
rect 33048 54606 33100 54612
rect 33508 54596 33560 54602
rect 33508 54538 33560 54544
rect 33140 54528 33192 54534
rect 33140 54470 33192 54476
rect 32772 54324 32824 54330
rect 32772 54266 32824 54272
rect 32404 54188 32456 54194
rect 32404 54130 32456 54136
rect 32036 53984 32088 53990
rect 32036 53926 32088 53932
rect 32784 53786 32812 54266
rect 32772 53780 32824 53786
rect 32772 53722 32824 53728
rect 33152 53582 33180 54470
rect 33520 54330 33548 54538
rect 33508 54324 33560 54330
rect 33508 54266 33560 54272
rect 33612 54262 33640 55014
rect 33704 54330 33732 55830
rect 33784 55752 33836 55758
rect 33784 55694 33836 55700
rect 33692 54324 33744 54330
rect 33692 54266 33744 54272
rect 33600 54256 33652 54262
rect 33600 54198 33652 54204
rect 33612 53786 33640 54198
rect 33600 53780 33652 53786
rect 33600 53722 33652 53728
rect 33140 53576 33192 53582
rect 33140 53518 33192 53524
rect 31944 53440 31996 53446
rect 31944 53382 31996 53388
rect 31956 53242 31984 53382
rect 30288 53236 30340 53242
rect 30288 53178 30340 53184
rect 31944 53236 31996 53242
rect 31944 53178 31996 53184
rect 33796 53174 33824 55694
rect 33968 55072 34020 55078
rect 33968 55014 34020 55020
rect 33980 54670 34008 55014
rect 33968 54664 34020 54670
rect 33968 54606 34020 54612
rect 34164 53514 34192 56306
rect 34336 56296 34388 56302
rect 34336 56238 34388 56244
rect 34348 55758 34376 56238
rect 34336 55752 34388 55758
rect 34336 55694 34388 55700
rect 34244 55344 34296 55350
rect 34244 55286 34296 55292
rect 34256 55214 34284 55286
rect 34244 55208 34296 55214
rect 34244 55150 34296 55156
rect 34256 54194 34284 55150
rect 34440 55146 34468 56306
rect 34520 55616 34572 55622
rect 34520 55558 34572 55564
rect 34532 55282 34560 55558
rect 34520 55276 34572 55282
rect 34520 55218 34572 55224
rect 34428 55140 34480 55146
rect 34428 55082 34480 55088
rect 34440 54670 34468 55082
rect 34532 54738 34560 55218
rect 34624 55128 34652 57190
rect 34702 57080 34758 57089
rect 34702 57015 34704 57024
rect 34756 57015 34758 57024
rect 34704 56986 34756 56992
rect 34704 56296 34756 56302
rect 34704 56238 34756 56244
rect 34716 56166 34744 56238
rect 34704 56160 34756 56166
rect 34704 56102 34756 56108
rect 34716 55758 34744 56102
rect 34704 55752 34756 55758
rect 34704 55694 34756 55700
rect 34808 55622 34836 57208
rect 35348 57190 35400 57196
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 35360 56438 35388 57190
rect 35348 56432 35400 56438
rect 35348 56374 35400 56380
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 35452 55962 35480 59200
rect 35532 57792 35584 57798
rect 35532 57734 35584 57740
rect 35716 57792 35768 57798
rect 35716 57734 35768 57740
rect 35544 56506 35572 57734
rect 35624 56908 35676 56914
rect 35624 56850 35676 56856
rect 35532 56500 35584 56506
rect 35532 56442 35584 56448
rect 35636 56370 35664 56850
rect 35624 56364 35676 56370
rect 35624 56306 35676 56312
rect 35728 56302 35756 57734
rect 35912 57390 35940 59200
rect 35992 57928 36044 57934
rect 35992 57870 36044 57876
rect 35808 57384 35860 57390
rect 35808 57326 35860 57332
rect 35900 57384 35952 57390
rect 35900 57326 35952 57332
rect 35820 56896 35848 57326
rect 35820 56868 35940 56896
rect 35808 56772 35860 56778
rect 35808 56714 35860 56720
rect 35820 56370 35848 56714
rect 35808 56364 35860 56370
rect 35808 56306 35860 56312
rect 35716 56296 35768 56302
rect 35716 56238 35768 56244
rect 35440 55956 35492 55962
rect 35440 55898 35492 55904
rect 35532 55820 35584 55826
rect 35728 55808 35756 56238
rect 35532 55762 35584 55768
rect 35636 55780 35756 55808
rect 34796 55616 34848 55622
rect 34796 55558 34848 55564
rect 35440 55344 35492 55350
rect 35544 55332 35572 55762
rect 35492 55304 35572 55332
rect 35440 55286 35492 55292
rect 34704 55140 34756 55146
rect 34624 55100 34704 55128
rect 34624 54738 34652 55100
rect 34704 55082 34756 55088
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34520 54732 34572 54738
rect 34520 54674 34572 54680
rect 34612 54732 34664 54738
rect 34612 54674 34664 54680
rect 34980 54732 35032 54738
rect 34980 54674 35032 54680
rect 34428 54664 34480 54670
rect 34428 54606 34480 54612
rect 34704 54664 34756 54670
rect 34704 54606 34756 54612
rect 34428 54528 34480 54534
rect 34428 54470 34480 54476
rect 34244 54188 34296 54194
rect 34244 54130 34296 54136
rect 34440 53786 34468 54470
rect 34716 54194 34744 54606
rect 34888 54596 34940 54602
rect 34888 54538 34940 54544
rect 34704 54188 34756 54194
rect 34704 54130 34756 54136
rect 34900 54126 34928 54538
rect 34992 54194 35020 54674
rect 35636 54194 35664 55780
rect 35716 55684 35768 55690
rect 35716 55626 35768 55632
rect 35728 55418 35756 55626
rect 35820 55418 35848 56306
rect 35716 55412 35768 55418
rect 35716 55354 35768 55360
rect 35808 55412 35860 55418
rect 35808 55354 35860 55360
rect 35912 54670 35940 56868
rect 36004 56846 36032 57870
rect 36176 57384 36228 57390
rect 36176 57326 36228 57332
rect 35992 56840 36044 56846
rect 35992 56782 36044 56788
rect 36004 56370 36032 56782
rect 36082 56400 36138 56409
rect 35992 56364 36044 56370
rect 36082 56335 36138 56344
rect 35992 56306 36044 56312
rect 36096 55826 36124 56335
rect 36084 55820 36136 55826
rect 36084 55762 36136 55768
rect 36084 55616 36136 55622
rect 36084 55558 36136 55564
rect 35990 55312 36046 55321
rect 35990 55247 36046 55256
rect 36004 55214 36032 55247
rect 35992 55208 36044 55214
rect 35992 55150 36044 55156
rect 35900 54664 35952 54670
rect 35900 54606 35952 54612
rect 34980 54188 35032 54194
rect 34980 54130 35032 54136
rect 35624 54188 35676 54194
rect 35624 54130 35676 54136
rect 34888 54120 34940 54126
rect 34888 54062 34940 54068
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 35636 53786 35664 54130
rect 35912 53786 35940 54606
rect 36096 54194 36124 55558
rect 36084 54188 36136 54194
rect 36084 54130 36136 54136
rect 34428 53780 34480 53786
rect 34428 53722 34480 53728
rect 35624 53780 35676 53786
rect 35624 53722 35676 53728
rect 35900 53780 35952 53786
rect 35900 53722 35952 53728
rect 34152 53508 34204 53514
rect 34152 53450 34204 53456
rect 35636 53242 35664 53722
rect 36084 53576 36136 53582
rect 36084 53518 36136 53524
rect 35624 53236 35676 53242
rect 35624 53178 35676 53184
rect 33784 53168 33836 53174
rect 33784 53110 33836 53116
rect 29460 53100 29512 53106
rect 29460 53042 29512 53048
rect 34520 53032 34572 53038
rect 34520 52974 34572 52980
rect 29368 52692 29420 52698
rect 29368 52634 29420 52640
rect 34532 16574 34560 52974
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 35636 52698 35664 53178
rect 36096 53106 36124 53518
rect 36084 53100 36136 53106
rect 36084 53042 36136 53048
rect 36188 52698 36216 57326
rect 36268 56976 36320 56982
rect 36268 56918 36320 56924
rect 36280 56846 36308 56918
rect 36268 56840 36320 56846
rect 36268 56782 36320 56788
rect 36280 55758 36308 56782
rect 36268 55752 36320 55758
rect 36268 55694 36320 55700
rect 36372 54194 36400 59200
rect 36832 57066 36860 59200
rect 37292 57390 37320 59200
rect 37556 57452 37608 57458
rect 37556 57394 37608 57400
rect 37280 57384 37332 57390
rect 37280 57326 37332 57332
rect 37280 57248 37332 57254
rect 37280 57190 37332 57196
rect 36728 57044 36780 57050
rect 36832 57038 36952 57066
rect 36728 56986 36780 56992
rect 36636 56840 36688 56846
rect 36740 56828 36768 56986
rect 36688 56800 36768 56828
rect 36636 56782 36688 56788
rect 36452 56364 36504 56370
rect 36452 56306 36504 56312
rect 36360 54188 36412 54194
rect 36360 54130 36412 54136
rect 36464 53174 36492 56306
rect 36544 55888 36596 55894
rect 36544 55830 36596 55836
rect 36556 54874 36584 55830
rect 36740 55622 36768 56800
rect 36820 56840 36872 56846
rect 36820 56782 36872 56788
rect 36832 56506 36860 56782
rect 36820 56500 36872 56506
rect 36820 56442 36872 56448
rect 36832 55758 36860 56442
rect 36924 55894 36952 57038
rect 37188 55956 37240 55962
rect 37188 55898 37240 55904
rect 36912 55888 36964 55894
rect 36912 55830 36964 55836
rect 36820 55752 36872 55758
rect 36820 55694 36872 55700
rect 36728 55616 36780 55622
rect 36728 55558 36780 55564
rect 37200 54874 37228 55898
rect 37292 55214 37320 57190
rect 37568 56846 37596 57394
rect 37556 56840 37608 56846
rect 37476 56800 37556 56828
rect 37476 56438 37504 56800
rect 37556 56782 37608 56788
rect 37464 56432 37516 56438
rect 37464 56374 37516 56380
rect 37372 56228 37424 56234
rect 37372 56170 37424 56176
rect 37384 55282 37412 56170
rect 37476 55962 37504 56374
rect 37554 55992 37610 56001
rect 37464 55956 37516 55962
rect 37554 55927 37610 55936
rect 37464 55898 37516 55904
rect 37372 55276 37424 55282
rect 37372 55218 37424 55224
rect 37280 55208 37332 55214
rect 37280 55150 37332 55156
rect 36544 54868 36596 54874
rect 36544 54810 36596 54816
rect 37188 54868 37240 54874
rect 37188 54810 37240 54816
rect 37384 54330 37412 55218
rect 37372 54324 37424 54330
rect 37372 54266 37424 54272
rect 37476 54262 37504 55898
rect 37568 55350 37596 55927
rect 37556 55344 37608 55350
rect 37556 55286 37608 55292
rect 37464 54256 37516 54262
rect 37464 54198 37516 54204
rect 37476 53718 37504 54198
rect 37752 53786 37780 59200
rect 38016 56840 38068 56846
rect 38016 56782 38068 56788
rect 38108 56840 38160 56846
rect 38108 56782 38160 56788
rect 37924 56364 37976 56370
rect 37924 56306 37976 56312
rect 37936 55418 37964 56306
rect 38028 55962 38056 56782
rect 38120 56234 38148 56782
rect 38212 56438 38240 59200
rect 38292 57384 38344 57390
rect 38292 57326 38344 57332
rect 38200 56432 38252 56438
rect 38200 56374 38252 56380
rect 38200 56296 38252 56302
rect 38200 56238 38252 56244
rect 38108 56228 38160 56234
rect 38108 56170 38160 56176
rect 38016 55956 38068 55962
rect 38016 55898 38068 55904
rect 37924 55412 37976 55418
rect 37924 55354 37976 55360
rect 38028 55282 38056 55898
rect 38212 55758 38240 56238
rect 38304 55962 38332 57326
rect 38672 56914 38700 59200
rect 38384 56908 38436 56914
rect 38384 56850 38436 56856
rect 38660 56908 38712 56914
rect 38660 56850 38712 56856
rect 38396 56001 38424 56850
rect 38382 55992 38438 56001
rect 38292 55956 38344 55962
rect 38382 55927 38438 55936
rect 38292 55898 38344 55904
rect 38200 55752 38252 55758
rect 38200 55694 38252 55700
rect 38016 55276 38068 55282
rect 38016 55218 38068 55224
rect 38212 54874 38240 55694
rect 38476 55684 38528 55690
rect 38476 55626 38528 55632
rect 38488 55418 38516 55626
rect 38476 55412 38528 55418
rect 38476 55354 38528 55360
rect 38200 54868 38252 54874
rect 38200 54810 38252 54816
rect 38568 54800 38620 54806
rect 38568 54742 38620 54748
rect 38384 54732 38436 54738
rect 38384 54674 38436 54680
rect 38396 54262 38424 54674
rect 38580 54262 38608 54742
rect 38384 54256 38436 54262
rect 38384 54198 38436 54204
rect 38568 54256 38620 54262
rect 38568 54198 38620 54204
rect 37740 53780 37792 53786
rect 37740 53722 37792 53728
rect 37464 53712 37516 53718
rect 37464 53654 37516 53660
rect 38672 53242 38700 56850
rect 38752 56840 38804 56846
rect 38752 56782 38804 56788
rect 39028 56840 39080 56846
rect 39028 56782 39080 56788
rect 38764 56302 38792 56782
rect 38844 56432 38896 56438
rect 38844 56374 38896 56380
rect 38752 56296 38804 56302
rect 38752 56238 38804 56244
rect 38752 55752 38804 55758
rect 38752 55694 38804 55700
rect 38764 55350 38792 55694
rect 38752 55344 38804 55350
rect 38752 55286 38804 55292
rect 38752 55208 38804 55214
rect 38752 55150 38804 55156
rect 38764 54602 38792 55150
rect 38752 54596 38804 54602
rect 38752 54538 38804 54544
rect 38856 53786 38884 56374
rect 39040 55622 39068 56782
rect 39132 56545 39160 59200
rect 39488 56704 39540 56710
rect 39488 56646 39540 56652
rect 39118 56536 39174 56545
rect 39500 56506 39528 56646
rect 39118 56471 39174 56480
rect 39488 56500 39540 56506
rect 39488 56442 39540 56448
rect 39212 55752 39264 55758
rect 39212 55694 39264 55700
rect 39028 55616 39080 55622
rect 39028 55558 39080 55564
rect 38936 55344 38988 55350
rect 38936 55286 38988 55292
rect 38948 54874 38976 55286
rect 39224 55282 39252 55694
rect 39304 55684 39356 55690
rect 39304 55626 39356 55632
rect 39212 55276 39264 55282
rect 39212 55218 39264 55224
rect 39120 55140 39172 55146
rect 39120 55082 39172 55088
rect 38936 54868 38988 54874
rect 38936 54810 38988 54816
rect 39132 54670 39160 55082
rect 39224 54670 39252 55218
rect 39316 55146 39344 55626
rect 39592 55282 39620 59200
rect 40052 59106 40080 59200
rect 40144 59106 40172 59214
rect 40052 59078 40172 59106
rect 40040 57860 40092 57866
rect 40040 57802 40092 57808
rect 40132 57860 40184 57866
rect 40132 57802 40184 57808
rect 40052 57594 40080 57802
rect 40040 57588 40092 57594
rect 40040 57530 40092 57536
rect 40144 57458 40172 57802
rect 40132 57452 40184 57458
rect 40132 57394 40184 57400
rect 39948 57384 40000 57390
rect 39948 57326 40000 57332
rect 39856 57044 39908 57050
rect 39856 56986 39908 56992
rect 39868 56846 39896 56986
rect 39856 56840 39908 56846
rect 39856 56782 39908 56788
rect 39672 55820 39724 55826
rect 39724 55780 39804 55808
rect 39672 55762 39724 55768
rect 39776 55622 39804 55780
rect 39764 55616 39816 55622
rect 39764 55558 39816 55564
rect 39580 55276 39632 55282
rect 39580 55218 39632 55224
rect 39304 55140 39356 55146
rect 39304 55082 39356 55088
rect 39580 55072 39632 55078
rect 39580 55014 39632 55020
rect 39592 54670 39620 55014
rect 39120 54664 39172 54670
rect 39120 54606 39172 54612
rect 39212 54664 39264 54670
rect 39212 54606 39264 54612
rect 39580 54664 39632 54670
rect 39580 54606 39632 54612
rect 39592 54330 39620 54606
rect 39776 54602 39804 55558
rect 39764 54596 39816 54602
rect 39764 54538 39816 54544
rect 39580 54324 39632 54330
rect 39580 54266 39632 54272
rect 39776 54210 39804 54538
rect 39684 54194 39804 54210
rect 39672 54188 39804 54194
rect 39724 54182 39804 54188
rect 39672 54130 39724 54136
rect 39868 53786 39896 56782
rect 39960 56370 39988 57326
rect 40132 57248 40184 57254
rect 40132 57190 40184 57196
rect 40144 56506 40172 57190
rect 40132 56500 40184 56506
rect 40132 56442 40184 56448
rect 39948 56364 40000 56370
rect 39948 56306 40000 56312
rect 40132 56364 40184 56370
rect 40132 56306 40184 56312
rect 39960 54262 39988 56306
rect 40040 55276 40092 55282
rect 40040 55218 40092 55224
rect 39948 54256 40000 54262
rect 39948 54198 40000 54204
rect 39960 53786 39988 54198
rect 40052 53990 40080 55218
rect 40144 54874 40172 56306
rect 40224 56296 40276 56302
rect 40224 56238 40276 56244
rect 40132 54868 40184 54874
rect 40132 54810 40184 54816
rect 40236 54126 40264 56238
rect 40328 54194 40356 59214
rect 40498 59200 40554 60000
rect 40958 59200 41014 60000
rect 41418 59200 41474 60000
rect 41878 59200 41934 60000
rect 42338 59200 42394 60000
rect 42798 59200 42854 60000
rect 43258 59200 43314 60000
rect 43718 59200 43774 60000
rect 44178 59200 44234 60000
rect 44638 59200 44694 60000
rect 45098 59200 45154 60000
rect 45558 59200 45614 60000
rect 46018 59200 46074 60000
rect 46478 59200 46534 60000
rect 46938 59200 46994 60000
rect 47398 59200 47454 60000
rect 47858 59200 47914 60000
rect 48318 59200 48374 60000
rect 48778 59200 48834 60000
rect 49238 59200 49294 60000
rect 49698 59200 49754 60000
rect 50158 59200 50214 60000
rect 50618 59200 50674 60000
rect 51078 59200 51134 60000
rect 51538 59200 51594 60000
rect 51998 59200 52054 60000
rect 52104 59214 52408 59242
rect 40408 57792 40460 57798
rect 40408 57734 40460 57740
rect 40420 57526 40448 57734
rect 40408 57520 40460 57526
rect 40408 57462 40460 57468
rect 40512 57474 40540 59200
rect 40512 57446 40632 57474
rect 40500 57384 40552 57390
rect 40500 57326 40552 57332
rect 40512 56506 40540 57326
rect 40500 56500 40552 56506
rect 40500 56442 40552 56448
rect 40604 56409 40632 57446
rect 40868 57452 40920 57458
rect 40972 57440 41000 59200
rect 41236 57452 41288 57458
rect 40972 57412 41092 57440
rect 40868 57394 40920 57400
rect 40776 56840 40828 56846
rect 40774 56808 40776 56817
rect 40828 56808 40830 56817
rect 40774 56743 40830 56752
rect 40880 56692 40908 57394
rect 40960 57316 41012 57322
rect 40960 57258 41012 57264
rect 40972 56846 41000 57258
rect 40960 56840 41012 56846
rect 40960 56782 41012 56788
rect 40960 56704 41012 56710
rect 40880 56664 40960 56692
rect 40960 56646 41012 56652
rect 40590 56400 40646 56409
rect 40590 56335 40646 56344
rect 40972 56166 41000 56646
rect 40408 56160 40460 56166
rect 40408 56102 40460 56108
rect 40960 56160 41012 56166
rect 41064 56137 41092 57412
rect 41236 57394 41288 57400
rect 41328 57452 41380 57458
rect 41328 57394 41380 57400
rect 41144 56976 41196 56982
rect 41142 56944 41144 56953
rect 41196 56944 41198 56953
rect 41248 56914 41276 57394
rect 41142 56879 41198 56888
rect 41236 56908 41288 56914
rect 41236 56850 41288 56856
rect 41144 56704 41196 56710
rect 41144 56646 41196 56652
rect 41156 56370 41184 56646
rect 41144 56364 41196 56370
rect 41144 56306 41196 56312
rect 40960 56102 41012 56108
rect 41050 56128 41106 56137
rect 40420 55078 40448 56102
rect 41050 56063 41106 56072
rect 40960 55956 41012 55962
rect 40960 55898 41012 55904
rect 40972 55758 41000 55898
rect 41340 55894 41368 57394
rect 41432 55978 41460 59200
rect 41788 57044 41840 57050
rect 41788 56986 41840 56992
rect 41800 56846 41828 56986
rect 41512 56840 41564 56846
rect 41512 56782 41564 56788
rect 41788 56840 41840 56846
rect 41788 56782 41840 56788
rect 41524 56302 41552 56782
rect 41892 56506 41920 59200
rect 42352 57866 42380 59200
rect 42340 57860 42392 57866
rect 42340 57802 42392 57808
rect 42812 57458 42840 59200
rect 42800 57452 42852 57458
rect 42800 57394 42852 57400
rect 43168 57316 43220 57322
rect 43168 57258 43220 57264
rect 42246 56944 42302 56953
rect 42246 56879 42302 56888
rect 41972 56840 42024 56846
rect 41970 56808 41972 56817
rect 42024 56808 42026 56817
rect 42260 56778 42288 56879
rect 43180 56846 43208 57258
rect 43168 56840 43220 56846
rect 43168 56782 43220 56788
rect 41970 56743 42026 56752
rect 42248 56772 42300 56778
rect 42248 56714 42300 56720
rect 41972 56704 42024 56710
rect 41972 56646 42024 56652
rect 41880 56500 41932 56506
rect 41880 56442 41932 56448
rect 41984 56370 42012 56646
rect 42892 56500 42944 56506
rect 42892 56442 42944 56448
rect 41972 56364 42024 56370
rect 41972 56306 42024 56312
rect 41512 56296 41564 56302
rect 41512 56238 41564 56244
rect 41878 56264 41934 56273
rect 41878 56199 41880 56208
rect 41932 56199 41934 56208
rect 42064 56228 42116 56234
rect 41880 56170 41932 56176
rect 42064 56170 42116 56176
rect 42800 56228 42852 56234
rect 42800 56170 42852 56176
rect 41432 55950 41552 55978
rect 41328 55888 41380 55894
rect 41328 55830 41380 55836
rect 41052 55820 41104 55826
rect 41052 55762 41104 55768
rect 40868 55752 40920 55758
rect 40868 55694 40920 55700
rect 40960 55752 41012 55758
rect 40960 55694 41012 55700
rect 40880 55418 40908 55694
rect 40960 55616 41012 55622
rect 40960 55558 41012 55564
rect 40868 55412 40920 55418
rect 40868 55354 40920 55360
rect 40408 55072 40460 55078
rect 40408 55014 40460 55020
rect 40420 54330 40448 55014
rect 40880 54738 40908 55354
rect 40868 54732 40920 54738
rect 40868 54674 40920 54680
rect 40972 54670 41000 55558
rect 41064 55078 41092 55762
rect 41524 55622 41552 55950
rect 41972 55752 42024 55758
rect 41972 55694 42024 55700
rect 41512 55616 41564 55622
rect 41512 55558 41564 55564
rect 41788 55412 41840 55418
rect 41788 55354 41840 55360
rect 41696 55208 41748 55214
rect 41696 55150 41748 55156
rect 41052 55072 41104 55078
rect 41052 55014 41104 55020
rect 40960 54664 41012 54670
rect 40960 54606 41012 54612
rect 40408 54324 40460 54330
rect 40408 54266 40460 54272
rect 41708 54194 41736 55150
rect 41800 54670 41828 55354
rect 41880 55072 41932 55078
rect 41880 55014 41932 55020
rect 41892 54670 41920 55014
rect 41984 54874 42012 55694
rect 42076 55282 42104 56170
rect 42248 56160 42300 56166
rect 42248 56102 42300 56108
rect 42708 56160 42760 56166
rect 42708 56102 42760 56108
rect 42064 55276 42116 55282
rect 42064 55218 42116 55224
rect 42076 55078 42104 55218
rect 42064 55072 42116 55078
rect 42064 55014 42116 55020
rect 41972 54868 42024 54874
rect 41972 54810 42024 54816
rect 41788 54664 41840 54670
rect 41788 54606 41840 54612
rect 41880 54664 41932 54670
rect 41880 54606 41932 54612
rect 41892 54330 41920 54606
rect 42076 54330 42104 55014
rect 42260 54534 42288 56102
rect 42432 55208 42484 55214
rect 42432 55150 42484 55156
rect 42248 54528 42300 54534
rect 42248 54470 42300 54476
rect 41880 54324 41932 54330
rect 41880 54266 41932 54272
rect 42064 54324 42116 54330
rect 42064 54266 42116 54272
rect 42444 54194 42472 55150
rect 42720 54330 42748 56102
rect 42812 54806 42840 56170
rect 42904 54874 42932 56442
rect 43180 55418 43208 56782
rect 43272 56234 43300 59200
rect 43352 57588 43404 57594
rect 43352 57530 43404 57536
rect 43364 56982 43392 57530
rect 43536 57452 43588 57458
rect 43536 57394 43588 57400
rect 43352 56976 43404 56982
rect 43352 56918 43404 56924
rect 43364 56846 43392 56918
rect 43352 56840 43404 56846
rect 43352 56782 43404 56788
rect 43352 56296 43404 56302
rect 43352 56238 43404 56244
rect 43260 56228 43312 56234
rect 43260 56170 43312 56176
rect 43260 55820 43312 55826
rect 43260 55762 43312 55768
rect 43168 55412 43220 55418
rect 43168 55354 43220 55360
rect 42892 54868 42944 54874
rect 42892 54810 42944 54816
rect 42800 54800 42852 54806
rect 42800 54742 42852 54748
rect 43180 54670 43208 55354
rect 43272 55078 43300 55762
rect 43364 55690 43392 56238
rect 43444 55752 43496 55758
rect 43444 55694 43496 55700
rect 43352 55684 43404 55690
rect 43352 55626 43404 55632
rect 43456 55282 43484 55694
rect 43444 55276 43496 55282
rect 43444 55218 43496 55224
rect 43260 55072 43312 55078
rect 43260 55014 43312 55020
rect 43548 54874 43576 57394
rect 43732 56982 43760 59200
rect 43996 57384 44048 57390
rect 43996 57326 44048 57332
rect 43904 57248 43956 57254
rect 43904 57190 43956 57196
rect 43720 56976 43772 56982
rect 43720 56918 43772 56924
rect 43916 56914 43944 57190
rect 43904 56908 43956 56914
rect 43904 56850 43956 56856
rect 43628 56840 43680 56846
rect 43628 56782 43680 56788
rect 43640 55894 43668 56782
rect 44008 56438 44036 57326
rect 44088 56840 44140 56846
rect 44086 56808 44088 56817
rect 44140 56808 44142 56817
rect 44086 56743 44142 56752
rect 43996 56432 44048 56438
rect 43996 56374 44048 56380
rect 44088 56364 44140 56370
rect 44088 56306 44140 56312
rect 44100 56273 44128 56306
rect 44086 56264 44142 56273
rect 44086 56199 44142 56208
rect 43628 55888 43680 55894
rect 43628 55830 43680 55836
rect 43640 55146 43668 55830
rect 44100 55826 44128 56199
rect 44088 55820 44140 55826
rect 44088 55762 44140 55768
rect 43720 55752 43772 55758
rect 43720 55694 43772 55700
rect 43732 55350 43760 55694
rect 43720 55344 43772 55350
rect 43720 55286 43772 55292
rect 44192 55282 44220 59200
rect 44456 57384 44508 57390
rect 44456 57326 44508 57332
rect 44272 57248 44324 57254
rect 44272 57190 44324 57196
rect 44284 57050 44312 57190
rect 44272 57044 44324 57050
rect 44272 56986 44324 56992
rect 44284 56506 44312 56986
rect 44468 56846 44496 57326
rect 44456 56840 44508 56846
rect 44456 56782 44508 56788
rect 44272 56500 44324 56506
rect 44272 56442 44324 56448
rect 44272 56296 44324 56302
rect 44468 56250 44496 56782
rect 44652 56302 44680 59200
rect 44732 57860 44784 57866
rect 44732 57802 44784 57808
rect 44324 56244 44496 56250
rect 44272 56238 44496 56244
rect 44640 56296 44692 56302
rect 44640 56238 44692 56244
rect 44284 56222 44496 56238
rect 44364 56160 44416 56166
rect 44364 56102 44416 56108
rect 44270 55992 44326 56001
rect 44270 55927 44272 55936
rect 44324 55927 44326 55936
rect 44272 55898 44324 55904
rect 44376 55826 44404 56102
rect 44364 55820 44416 55826
rect 44364 55762 44416 55768
rect 44468 55690 44496 56222
rect 44548 56160 44600 56166
rect 44548 56102 44600 56108
rect 44560 55758 44588 56102
rect 44744 55962 44772 57802
rect 44916 57452 44968 57458
rect 44916 57394 44968 57400
rect 44824 57248 44876 57254
rect 44824 57190 44876 57196
rect 44836 56545 44864 57190
rect 44822 56536 44878 56545
rect 44822 56471 44878 56480
rect 44732 55956 44784 55962
rect 44732 55898 44784 55904
rect 44548 55752 44600 55758
rect 44548 55694 44600 55700
rect 44456 55684 44508 55690
rect 44456 55626 44508 55632
rect 44180 55276 44232 55282
rect 44180 55218 44232 55224
rect 43628 55140 43680 55146
rect 43628 55082 43680 55088
rect 44928 55078 44956 57394
rect 45008 56772 45060 56778
rect 45008 56714 45060 56720
rect 45020 56506 45048 56714
rect 45008 56500 45060 56506
rect 45008 56442 45060 56448
rect 45020 56370 45048 56442
rect 45008 56364 45060 56370
rect 45008 56306 45060 56312
rect 45112 55962 45140 59200
rect 45572 57458 45600 59200
rect 45560 57452 45612 57458
rect 45560 57394 45612 57400
rect 45928 57248 45980 57254
rect 45928 57190 45980 57196
rect 45192 56840 45244 56846
rect 45192 56782 45244 56788
rect 45836 56840 45888 56846
rect 45836 56782 45888 56788
rect 45204 56409 45232 56782
rect 45190 56400 45246 56409
rect 45190 56335 45246 56344
rect 45284 56364 45336 56370
rect 45284 56306 45336 56312
rect 45100 55956 45152 55962
rect 45100 55898 45152 55904
rect 45296 55826 45324 56306
rect 45848 56137 45876 56782
rect 45834 56128 45890 56137
rect 45834 56063 45890 56072
rect 45284 55820 45336 55826
rect 45284 55762 45336 55768
rect 45296 55418 45324 55762
rect 45284 55412 45336 55418
rect 45284 55354 45336 55360
rect 45940 55214 45968 57190
rect 46032 57050 46060 59200
rect 46388 57452 46440 57458
rect 46388 57394 46440 57400
rect 46400 57322 46428 57394
rect 46388 57316 46440 57322
rect 46388 57258 46440 57264
rect 46020 57044 46072 57050
rect 46020 56986 46072 56992
rect 46492 56370 46520 59200
rect 46952 57458 46980 59200
rect 46756 57452 46808 57458
rect 46756 57394 46808 57400
rect 46940 57452 46992 57458
rect 46940 57394 46992 57400
rect 46480 56364 46532 56370
rect 46480 56306 46532 56312
rect 46768 55622 46796 57394
rect 47412 56370 47440 59200
rect 47584 57452 47636 57458
rect 47584 57394 47636 57400
rect 47400 56364 47452 56370
rect 47400 56306 47452 56312
rect 47596 55962 47624 57394
rect 47872 57050 47900 59200
rect 47860 57044 47912 57050
rect 47860 56986 47912 56992
rect 48332 56914 48360 59200
rect 48320 56908 48372 56914
rect 48320 56850 48372 56856
rect 48332 55962 48360 56850
rect 48688 56840 48740 56846
rect 48688 56782 48740 56788
rect 48700 56273 48728 56782
rect 48792 56370 48820 59200
rect 49148 57792 49200 57798
rect 49148 57734 49200 57740
rect 49160 57322 49188 57734
rect 49148 57316 49200 57322
rect 49148 57258 49200 57264
rect 49252 56370 49280 59200
rect 49712 57458 49740 59200
rect 49700 57452 49752 57458
rect 49700 57394 49752 57400
rect 49712 56506 49740 57394
rect 50172 57050 50200 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 50160 57044 50212 57050
rect 50160 56986 50212 56992
rect 50632 56982 50660 59200
rect 51092 57458 51120 59200
rect 51080 57452 51132 57458
rect 51080 57394 51132 57400
rect 51448 57452 51500 57458
rect 51448 57394 51500 57400
rect 50620 56976 50672 56982
rect 50620 56918 50672 56924
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 51460 56506 51488 57394
rect 51552 57050 51580 59200
rect 52012 59106 52040 59200
rect 52104 59106 52132 59214
rect 52012 59078 52132 59106
rect 51540 57044 51592 57050
rect 52380 57032 52408 59214
rect 52458 59200 52514 60000
rect 52918 59200 52974 60000
rect 53378 59200 53434 60000
rect 53838 59200 53894 60000
rect 54298 59200 54354 60000
rect 54758 59200 54814 60000
rect 55218 59200 55274 60000
rect 55678 59200 55734 60000
rect 56138 59200 56194 60000
rect 52472 57526 52500 59200
rect 52460 57520 52512 57526
rect 52460 57462 52512 57468
rect 52828 57520 52880 57526
rect 52828 57462 52880 57468
rect 52460 57044 52512 57050
rect 52380 57004 52460 57032
rect 51540 56986 51592 56992
rect 52460 56986 52512 56992
rect 52840 56506 52868 57462
rect 52932 57050 52960 59200
rect 52920 57044 52972 57050
rect 53392 57032 53420 59200
rect 53852 57458 53880 59200
rect 54312 57458 54340 59200
rect 53840 57452 53892 57458
rect 53840 57394 53892 57400
rect 54300 57452 54352 57458
rect 54300 57394 54352 57400
rect 53472 57044 53524 57050
rect 53392 57004 53472 57032
rect 52920 56986 52972 56992
rect 53472 56986 53524 56992
rect 53852 56506 53880 57394
rect 54116 57248 54168 57254
rect 54116 57190 54168 57196
rect 54208 57248 54260 57254
rect 54208 57190 54260 57196
rect 54128 56778 54156 57190
rect 54116 56772 54168 56778
rect 54116 56714 54168 56720
rect 49700 56500 49752 56506
rect 49700 56442 49752 56448
rect 51448 56500 51500 56506
rect 51448 56442 51500 56448
rect 52828 56500 52880 56506
rect 52828 56442 52880 56448
rect 53840 56500 53892 56506
rect 53840 56442 53892 56448
rect 48780 56364 48832 56370
rect 48780 56306 48832 56312
rect 49240 56364 49292 56370
rect 49240 56306 49292 56312
rect 48686 56264 48742 56273
rect 48686 56199 48742 56208
rect 47584 55956 47636 55962
rect 47584 55898 47636 55904
rect 48320 55956 48372 55962
rect 48320 55898 48372 55904
rect 46756 55616 46808 55622
rect 46756 55558 46808 55564
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 54220 55418 54248 57190
rect 54772 57050 54800 59200
rect 55232 57458 55260 59200
rect 55692 57458 55720 59200
rect 55220 57452 55272 57458
rect 55220 57394 55272 57400
rect 55680 57452 55732 57458
rect 55680 57394 55732 57400
rect 55232 57050 55260 57394
rect 56152 57050 56180 59200
rect 54760 57044 54812 57050
rect 54760 56986 54812 56992
rect 55220 57044 55272 57050
rect 55220 56986 55272 56992
rect 56140 57044 56192 57050
rect 56140 56986 56192 56992
rect 54208 55412 54260 55418
rect 54208 55354 54260 55360
rect 45928 55208 45980 55214
rect 45928 55150 45980 55156
rect 44916 55072 44968 55078
rect 44916 55014 44968 55020
rect 43536 54868 43588 54874
rect 43536 54810 43588 54816
rect 43168 54664 43220 54670
rect 43168 54606 43220 54612
rect 44928 54602 44956 55014
rect 44916 54596 44968 54602
rect 44916 54538 44968 54544
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 42708 54324 42760 54330
rect 42708 54266 42760 54272
rect 40316 54188 40368 54194
rect 40316 54130 40368 54136
rect 40776 54188 40828 54194
rect 40776 54130 40828 54136
rect 41696 54188 41748 54194
rect 41696 54130 41748 54136
rect 42432 54188 42484 54194
rect 42432 54130 42484 54136
rect 40224 54120 40276 54126
rect 40224 54062 40276 54068
rect 40040 53984 40092 53990
rect 40040 53926 40092 53932
rect 40788 53786 40816 54130
rect 42720 53786 42748 54266
rect 38844 53780 38896 53786
rect 38844 53722 38896 53728
rect 39856 53780 39908 53786
rect 39856 53722 39908 53728
rect 39948 53780 40000 53786
rect 39948 53722 40000 53728
rect 40776 53780 40828 53786
rect 40776 53722 40828 53728
rect 42708 53780 42760 53786
rect 42708 53722 42760 53728
rect 39960 53582 39988 53722
rect 39948 53576 40000 53582
rect 39948 53518 40000 53524
rect 39960 53242 39988 53518
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 38660 53236 38712 53242
rect 38660 53178 38712 53184
rect 39948 53236 40000 53242
rect 39948 53178 40000 53184
rect 36452 53168 36504 53174
rect 36452 53110 36504 53116
rect 35624 52692 35676 52698
rect 35624 52634 35676 52640
rect 36176 52692 36228 52698
rect 36176 52634 36228 52640
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34532 16546 34652 16574
rect 26424 8084 26476 8090
rect 26424 8026 26476 8032
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 24952 7472 25004 7478
rect 24952 7414 25004 7420
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 7668 800 7696 2790
rect 8220 800 8248 2790
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 8588 800 8616 2518
rect 8956 800 8984 2790
rect 9324 800 9352 3470
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9692 800 9720 2382
rect 9968 800 9996 2790
rect 10244 800 10272 3470
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 10520 800 10548 2790
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10796 800 10824 2450
rect 11072 800 11100 2790
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11348 800 11376 2382
rect 11624 800 11652 2790
rect 11900 800 11928 3470
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 12176 800 12204 2790
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12452 800 12480 2518
rect 12728 800 12756 3470
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 13004 800 13032 2790
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13280 800 13308 2382
rect 13556 800 13584 3470
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 13832 800 13860 2790
rect 14108 800 14136 2790
rect 14384 800 14412 3470
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 14660 800 14688 2450
rect 14936 800 14964 3470
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15212 800 15240 2790
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15488 800 15516 2382
rect 15764 800 15792 3470
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 16040 800 16068 2926
rect 16316 800 16344 3878
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16592 800 16620 2790
rect 16868 800 16896 3470
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 17144 800 17172 2450
rect 17328 800 17356 2790
rect 17604 800 17632 3878
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 17880 800 17908 3470
rect 18156 800 18184 3470
rect 18432 800 18460 3878
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 18696 2576 18748 2582
rect 18696 2518 18748 2524
rect 18708 800 18736 2518
rect 18984 800 19012 2926
rect 19352 2802 19380 4558
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19260 2774 19380 2802
rect 19260 800 19288 2774
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 19352 1442 19380 2246
rect 19444 1986 19472 3878
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 19996 2922 20024 3062
rect 19524 2916 19576 2922
rect 19524 2858 19576 2864
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 19536 2310 19564 2858
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19524 2304 19576 2310
rect 19524 2246 19576 2252
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 2106 20024 2382
rect 19984 2100 20036 2106
rect 19984 2042 20036 2048
rect 19444 1958 19840 1986
rect 19352 1414 19564 1442
rect 19536 800 19564 1414
rect 19812 800 19840 1958
rect 20088 800 20116 3538
rect 20364 800 20392 4558
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20640 800 20668 4014
rect 21456 3664 21508 3670
rect 21456 3606 21508 3612
rect 21180 3052 21232 3058
rect 21180 2994 21232 3000
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 20916 800 20944 2450
rect 21192 800 21220 2994
rect 21468 800 21496 3606
rect 21744 800 21772 4558
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 22020 800 22048 3946
rect 22204 3058 22232 4558
rect 22296 4146 22324 5102
rect 22572 4826 22600 7278
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 23940 6112 23992 6118
rect 23940 6054 23992 6060
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 22836 5024 22888 5030
rect 22836 4966 22888 4972
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22744 4072 22796 4078
rect 22744 4014 22796 4020
rect 22756 3738 22784 4014
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 22572 3058 22600 3470
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22204 2310 22232 2994
rect 22560 2916 22612 2922
rect 22560 2858 22612 2864
rect 22284 2372 22336 2378
rect 22284 2314 22336 2320
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22296 800 22324 2314
rect 22572 800 22600 2858
rect 22848 800 22876 4966
rect 22928 4072 22980 4078
rect 22928 4014 22980 4020
rect 22940 2650 22968 4014
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 23124 800 23152 5646
rect 23388 4752 23440 4758
rect 23388 4694 23440 4700
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23308 2310 23336 2382
rect 23296 2304 23348 2310
rect 23296 2246 23348 2252
rect 23400 800 23428 4694
rect 23848 3460 23900 3466
rect 23848 3402 23900 3408
rect 23664 3392 23716 3398
rect 23664 3334 23716 3340
rect 23676 800 23704 3334
rect 23860 2650 23888 3402
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 23952 800 23980 6054
rect 24504 5710 24532 6258
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24688 5778 24716 6054
rect 24872 5778 24900 6598
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 24492 5704 24544 5710
rect 24492 5646 24544 5652
rect 24124 5568 24176 5574
rect 24124 5510 24176 5516
rect 24136 5302 24164 5510
rect 24124 5296 24176 5302
rect 24124 5238 24176 5244
rect 24504 5234 24532 5646
rect 24492 5228 24544 5234
rect 24492 5170 24544 5176
rect 24504 4690 24532 5170
rect 24492 4684 24544 4690
rect 24492 4626 24544 4632
rect 24492 3936 24544 3942
rect 24492 3878 24544 3884
rect 24216 3120 24268 3126
rect 24216 3062 24268 3068
rect 24228 800 24256 3062
rect 24504 800 24532 3878
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24596 3058 24624 3470
rect 24964 3194 24992 7414
rect 26436 6914 26464 8026
rect 30288 7404 30340 7410
rect 30288 7346 30340 7352
rect 26792 7336 26844 7342
rect 26792 7278 26844 7284
rect 26700 7200 26752 7206
rect 26700 7142 26752 7148
rect 26436 6886 26556 6914
rect 25596 6860 25648 6866
rect 25596 6802 25648 6808
rect 25412 5160 25464 5166
rect 25412 5102 25464 5108
rect 24952 3188 25004 3194
rect 24952 3130 25004 3136
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 25228 2984 25280 2990
rect 25228 2926 25280 2932
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 24768 2100 24820 2106
rect 24768 2042 24820 2048
rect 24780 800 24808 2042
rect 25056 800 25084 2790
rect 25240 2650 25268 2926
rect 25424 2854 25452 5102
rect 25608 4146 25636 6802
rect 26528 6730 26556 6886
rect 26608 6792 26660 6798
rect 26608 6734 26660 6740
rect 26516 6724 26568 6730
rect 26516 6666 26568 6672
rect 26240 6248 26292 6254
rect 26240 6190 26292 6196
rect 26148 5772 26200 5778
rect 26148 5714 26200 5720
rect 26056 5704 26108 5710
rect 26056 5646 26108 5652
rect 26068 5234 26096 5646
rect 26056 5228 26108 5234
rect 26056 5170 26108 5176
rect 25596 4140 25648 4146
rect 25596 4082 25648 4088
rect 25412 2848 25464 2854
rect 25412 2790 25464 2796
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 25596 2576 25648 2582
rect 25596 2518 25648 2524
rect 25320 2304 25372 2310
rect 25320 2246 25372 2252
rect 25332 800 25360 2246
rect 25608 800 25636 2518
rect 25872 2508 25924 2514
rect 25872 2450 25924 2456
rect 25884 800 25912 2450
rect 26160 800 26188 5714
rect 26252 4146 26280 6190
rect 26528 5710 26556 6666
rect 26620 6322 26648 6734
rect 26608 6316 26660 6322
rect 26608 6258 26660 6264
rect 26516 5704 26568 5710
rect 26516 5646 26568 5652
rect 26712 5234 26740 7142
rect 26700 5228 26752 5234
rect 26700 5170 26752 5176
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 26516 3528 26568 3534
rect 26804 3482 26832 7278
rect 29736 7200 29788 7206
rect 29736 7142 29788 7148
rect 28632 6860 28684 6866
rect 28632 6802 28684 6808
rect 28172 6724 28224 6730
rect 28172 6666 28224 6672
rect 26884 6656 26936 6662
rect 26884 6598 26936 6604
rect 26896 5302 26924 6598
rect 27896 6248 27948 6254
rect 27896 6190 27948 6196
rect 27528 5704 27580 5710
rect 27528 5646 27580 5652
rect 26976 5636 27028 5642
rect 26976 5578 27028 5584
rect 26988 5370 27016 5578
rect 26976 5364 27028 5370
rect 26976 5306 27028 5312
rect 26884 5296 26936 5302
rect 26884 5238 26936 5244
rect 27540 4826 27568 5646
rect 27528 4820 27580 4826
rect 27528 4762 27580 4768
rect 27528 4548 27580 4554
rect 27528 4490 27580 4496
rect 27436 4072 27488 4078
rect 27436 4014 27488 4020
rect 27252 3936 27304 3942
rect 27252 3878 27304 3884
rect 26976 3664 27028 3670
rect 26976 3606 27028 3612
rect 26516 3470 26568 3476
rect 26332 3460 26384 3466
rect 26332 3402 26384 3408
rect 26344 2650 26372 3402
rect 26528 3058 26556 3470
rect 26712 3454 26832 3482
rect 26516 3052 26568 3058
rect 26516 2994 26568 3000
rect 26424 2848 26476 2854
rect 26424 2790 26476 2796
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 26436 800 26464 2790
rect 26712 800 26740 3454
rect 26988 800 27016 3606
rect 27264 800 27292 3878
rect 27448 3738 27476 4014
rect 27436 3732 27488 3738
rect 27436 3674 27488 3680
rect 27436 3528 27488 3534
rect 27436 3470 27488 3476
rect 27448 2446 27476 3470
rect 27436 2440 27488 2446
rect 27436 2382 27488 2388
rect 27540 800 27568 4490
rect 27804 2984 27856 2990
rect 27804 2926 27856 2932
rect 27816 2650 27844 2926
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 27908 2530 27936 6190
rect 28080 5772 28132 5778
rect 28080 5714 28132 5720
rect 27988 4004 28040 4010
rect 27988 3946 28040 3952
rect 28000 3738 28028 3946
rect 27988 3732 28040 3738
rect 27988 3674 28040 3680
rect 27816 2502 27936 2530
rect 27816 800 27844 2502
rect 28092 800 28120 5714
rect 28184 2378 28212 6666
rect 28356 5160 28408 5166
rect 28356 5102 28408 5108
rect 28172 2372 28224 2378
rect 28172 2314 28224 2320
rect 28368 800 28396 5102
rect 28644 800 28672 6802
rect 29552 6792 29604 6798
rect 29552 6734 29604 6740
rect 29564 6322 29592 6734
rect 29748 6390 29776 7142
rect 29736 6384 29788 6390
rect 29736 6326 29788 6332
rect 29552 6316 29604 6322
rect 29552 6258 29604 6264
rect 30300 6254 30328 7346
rect 30380 7200 30432 7206
rect 30380 7142 30432 7148
rect 30392 6662 30420 7142
rect 31024 6792 31076 6798
rect 31024 6734 31076 6740
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 30380 6656 30432 6662
rect 30380 6598 30432 6604
rect 30196 6248 30248 6254
rect 30196 6190 30248 6196
rect 30288 6248 30340 6254
rect 30288 6190 30340 6196
rect 30104 5772 30156 5778
rect 30104 5714 30156 5720
rect 30012 4684 30064 4690
rect 30012 4626 30064 4632
rect 29460 4548 29512 4554
rect 29460 4490 29512 4496
rect 29184 3664 29236 3670
rect 29184 3606 29236 3612
rect 29092 3460 29144 3466
rect 29092 3402 29144 3408
rect 28908 2916 28960 2922
rect 28908 2858 28960 2864
rect 28920 800 28948 2858
rect 29104 2650 29132 3402
rect 29092 2644 29144 2650
rect 29092 2586 29144 2592
rect 29196 800 29224 3606
rect 29472 3194 29500 4490
rect 29552 4140 29604 4146
rect 29552 4082 29604 4088
rect 29460 3188 29512 3194
rect 29460 3130 29512 3136
rect 29564 3058 29592 4082
rect 29736 4072 29788 4078
rect 29736 4014 29788 4020
rect 29644 3596 29696 3602
rect 29644 3538 29696 3544
rect 29552 3052 29604 3058
rect 29552 2994 29604 3000
rect 29460 2984 29512 2990
rect 29460 2926 29512 2932
rect 29472 800 29500 2926
rect 29564 2446 29592 2994
rect 29656 2650 29684 3538
rect 29644 2644 29696 2650
rect 29644 2586 29696 2592
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 29748 800 29776 4014
rect 30024 800 30052 4626
rect 30116 4146 30144 5714
rect 30104 4140 30156 4146
rect 30104 4082 30156 4088
rect 30208 3210 30236 6190
rect 30300 5778 30328 6190
rect 30288 5772 30340 5778
rect 30288 5714 30340 5720
rect 30392 5710 30420 6598
rect 31036 5778 31064 6734
rect 31208 6112 31260 6118
rect 31208 6054 31260 6060
rect 31220 5778 31248 6054
rect 31024 5772 31076 5778
rect 31024 5714 31076 5720
rect 31208 5772 31260 5778
rect 31208 5714 31260 5720
rect 31668 5772 31720 5778
rect 31668 5714 31720 5720
rect 30380 5704 30432 5710
rect 30380 5646 30432 5652
rect 31024 5636 31076 5642
rect 31024 5578 31076 5584
rect 30288 5160 30340 5166
rect 30288 5102 30340 5108
rect 30564 5160 30616 5166
rect 30564 5102 30616 5108
rect 30300 4282 30328 5102
rect 30288 4276 30340 4282
rect 30288 4218 30340 4224
rect 30208 3182 30328 3210
rect 30300 800 30328 3182
rect 30380 2916 30432 2922
rect 30380 2858 30432 2864
rect 30392 2650 30420 2858
rect 30380 2644 30432 2650
rect 30380 2586 30432 2592
rect 30576 800 30604 5102
rect 31036 5030 31064 5578
rect 31024 5024 31076 5030
rect 31024 4966 31076 4972
rect 31036 4622 31064 4966
rect 31024 4616 31076 4622
rect 31024 4558 31076 4564
rect 30656 4072 30708 4078
rect 30656 4014 30708 4020
rect 31392 4072 31444 4078
rect 31392 4014 31444 4020
rect 30668 3738 30696 4014
rect 30656 3732 30708 3738
rect 30656 3674 30708 3680
rect 31024 3460 31076 3466
rect 31024 3402 31076 3408
rect 30840 2916 30892 2922
rect 30840 2858 30892 2864
rect 30852 800 30880 2858
rect 31036 1714 31064 3402
rect 31116 2984 31168 2990
rect 31116 2926 31168 2932
rect 31128 2650 31156 2926
rect 31116 2644 31168 2650
rect 31116 2586 31168 2592
rect 31036 1686 31156 1714
rect 31128 800 31156 1686
rect 31404 800 31432 4014
rect 31680 800 31708 5714
rect 31772 5642 31800 6734
rect 32220 6656 32272 6662
rect 32220 6598 32272 6604
rect 31760 5636 31812 5642
rect 31760 5578 31812 5584
rect 31772 4690 31800 5578
rect 32232 4690 32260 6598
rect 34428 6248 34480 6254
rect 34428 6190 34480 6196
rect 33048 6112 33100 6118
rect 33048 6054 33100 6060
rect 31760 4684 31812 4690
rect 31760 4626 31812 4632
rect 32220 4684 32272 4690
rect 32220 4626 32272 4632
rect 32772 4684 32824 4690
rect 32772 4626 32824 4632
rect 32220 3664 32272 3670
rect 32220 3606 32272 3612
rect 31944 2984 31996 2990
rect 31944 2926 31996 2932
rect 31956 800 31984 2926
rect 32232 800 32260 3606
rect 32496 3596 32548 3602
rect 32496 3538 32548 3544
rect 32508 800 32536 3538
rect 32784 800 32812 4626
rect 33060 4146 33088 6054
rect 33140 5704 33192 5710
rect 33140 5646 33192 5652
rect 33152 4758 33180 5646
rect 33232 5568 33284 5574
rect 33232 5510 33284 5516
rect 33140 4752 33192 4758
rect 33140 4694 33192 4700
rect 33048 4140 33100 4146
rect 33048 4082 33100 4088
rect 33244 4078 33272 5510
rect 33324 5160 33376 5166
rect 33324 5102 33376 5108
rect 33232 4072 33284 4078
rect 33232 4014 33284 4020
rect 33048 4004 33100 4010
rect 33048 3946 33100 3952
rect 33060 800 33088 3946
rect 33336 800 33364 5102
rect 34152 4004 34204 4010
rect 34152 3946 34204 3952
rect 33876 3936 33928 3942
rect 33876 3878 33928 3884
rect 33692 3528 33744 3534
rect 33692 3470 33744 3476
rect 33600 2848 33652 2854
rect 33600 2790 33652 2796
rect 33612 800 33640 2790
rect 33704 2650 33732 3470
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 33888 800 33916 3878
rect 34164 800 34192 3946
rect 34336 3528 34388 3534
rect 34336 3470 34388 3476
rect 34348 2446 34376 3470
rect 34336 2440 34388 2446
rect 34336 2382 34388 2388
rect 34440 800 34468 6190
rect 34520 2916 34572 2922
rect 34520 2858 34572 2864
rect 34532 2582 34560 2858
rect 34520 2576 34572 2582
rect 34520 2518 34572 2524
rect 34624 2530 34652 16546
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 38200 6384 38252 6390
rect 38200 6326 38252 6332
rect 37924 6248 37976 6254
rect 37924 6190 37976 6196
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35348 5704 35400 5710
rect 35348 5646 35400 5652
rect 34796 5568 34848 5574
rect 34796 5510 34848 5516
rect 34808 5302 34836 5510
rect 34796 5296 34848 5302
rect 34796 5238 34848 5244
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34980 4548 35032 4554
rect 34980 4490 35032 4496
rect 34992 3942 35020 4490
rect 35360 4146 35388 5646
rect 35900 5024 35952 5030
rect 35900 4966 35952 4972
rect 35348 4140 35400 4146
rect 35348 4082 35400 4088
rect 34980 3936 35032 3942
rect 34980 3878 35032 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35360 3602 35388 4082
rect 35440 3936 35492 3942
rect 35440 3878 35492 3884
rect 35348 3596 35400 3602
rect 35348 3538 35400 3544
rect 34980 3528 35032 3534
rect 34980 3470 35032 3476
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 34704 2984 34756 2990
rect 34704 2926 34756 2932
rect 34716 2650 34744 2926
rect 34704 2644 34756 2650
rect 34704 2586 34756 2592
rect 34624 2502 34744 2530
rect 34716 800 34744 2502
rect 34808 1714 34836 3334
rect 34992 3058 35020 3470
rect 35348 3460 35400 3466
rect 35348 3402 35400 3408
rect 34980 3052 35032 3058
rect 34980 2994 35032 3000
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 2650 35388 3402
rect 35452 3126 35480 3878
rect 35532 3596 35584 3602
rect 35532 3538 35584 3544
rect 35440 3120 35492 3126
rect 35440 3062 35492 3068
rect 35440 2848 35492 2854
rect 35440 2790 35492 2796
rect 35348 2644 35400 2650
rect 35348 2586 35400 2592
rect 34808 1686 35020 1714
rect 34992 800 35020 1686
rect 35452 1442 35480 2790
rect 35268 1414 35480 1442
rect 35268 800 35296 1414
rect 35544 800 35572 3538
rect 35808 2916 35860 2922
rect 35808 2858 35860 2864
rect 35820 800 35848 2858
rect 35912 2854 35940 4966
rect 37280 4752 37332 4758
rect 37280 4694 37332 4700
rect 36820 4616 36872 4622
rect 36820 4558 36872 4564
rect 36832 4146 36860 4558
rect 36820 4140 36872 4146
rect 36820 4082 36872 4088
rect 37004 4072 37056 4078
rect 37004 4014 37056 4020
rect 37188 4072 37240 4078
rect 37188 4014 37240 4020
rect 36636 3664 36688 3670
rect 36636 3606 36688 3612
rect 36360 3188 36412 3194
rect 36360 3130 36412 3136
rect 35900 2848 35952 2854
rect 35900 2790 35952 2796
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 36096 800 36124 2314
rect 36372 800 36400 3130
rect 36648 800 36676 3606
rect 36912 3460 36964 3466
rect 36912 3402 36964 3408
rect 36924 800 36952 3402
rect 37016 2650 37044 4014
rect 37004 2644 37056 2650
rect 37004 2586 37056 2592
rect 37200 2582 37228 4014
rect 37188 2576 37240 2582
rect 37188 2518 37240 2524
rect 37292 2394 37320 4694
rect 37464 4616 37516 4622
rect 37464 4558 37516 4564
rect 37372 4548 37424 4554
rect 37372 4490 37424 4496
rect 37384 3738 37412 4490
rect 37372 3732 37424 3738
rect 37372 3674 37424 3680
rect 37372 3528 37424 3534
rect 37372 3470 37424 3476
rect 37384 2446 37412 3470
rect 37476 3194 37504 4558
rect 37740 3936 37792 3942
rect 37740 3878 37792 3884
rect 37464 3188 37516 3194
rect 37464 3130 37516 3136
rect 37556 3120 37608 3126
rect 37556 3062 37608 3068
rect 37200 2366 37320 2394
rect 37372 2440 37424 2446
rect 37372 2382 37424 2388
rect 37200 800 37228 2366
rect 37568 1850 37596 3062
rect 37476 1822 37596 1850
rect 37476 800 37504 1822
rect 37752 800 37780 3878
rect 37936 3738 37964 6190
rect 37924 3732 37976 3738
rect 37924 3674 37976 3680
rect 38108 3732 38160 3738
rect 38108 3674 38160 3680
rect 38120 3126 38148 3674
rect 38108 3120 38160 3126
rect 38108 3062 38160 3068
rect 38016 2916 38068 2922
rect 38016 2858 38068 2864
rect 38028 800 38056 2858
rect 38212 2650 38240 6326
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 38936 4616 38988 4622
rect 38936 4558 38988 4564
rect 38568 3596 38620 3602
rect 38568 3538 38620 3544
rect 38384 3052 38436 3058
rect 38384 2994 38436 3000
rect 38200 2644 38252 2650
rect 38200 2586 38252 2592
rect 38396 1442 38424 2994
rect 38304 1414 38424 1442
rect 38304 800 38332 1414
rect 38580 800 38608 3538
rect 38752 3392 38804 3398
rect 38752 3334 38804 3340
rect 38764 2650 38792 3334
rect 38948 2922 38976 4558
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 39120 4004 39172 4010
rect 39120 3946 39172 3952
rect 39028 3460 39080 3466
rect 39028 3402 39080 3408
rect 39040 2922 39068 3402
rect 38936 2916 38988 2922
rect 38936 2858 38988 2864
rect 39028 2916 39080 2922
rect 39028 2858 39080 2864
rect 38752 2644 38804 2650
rect 38752 2586 38804 2592
rect 38844 2508 38896 2514
rect 38844 2450 38896 2456
rect 38856 800 38884 2450
rect 39132 800 39160 3946
rect 40224 3936 40276 3942
rect 40224 3878 40276 3884
rect 39396 3664 39448 3670
rect 39396 3606 39448 3612
rect 39408 800 39436 3606
rect 40040 3392 40092 3398
rect 40040 3334 40092 3340
rect 39672 2984 39724 2990
rect 39672 2926 39724 2932
rect 39684 800 39712 2926
rect 40052 2650 40080 3334
rect 40040 2644 40092 2650
rect 40040 2586 40092 2592
rect 39948 2576 40000 2582
rect 39948 2518 40000 2524
rect 39960 800 39988 2518
rect 40236 800 40264 3878
rect 42156 3664 42208 3670
rect 42156 3606 42208 3612
rect 43260 3664 43312 3670
rect 43260 3606 43312 3612
rect 45468 3664 45520 3670
rect 45468 3606 45520 3612
rect 40776 3596 40828 3602
rect 40776 3538 40828 3544
rect 40500 2916 40552 2922
rect 40500 2858 40552 2864
rect 40512 800 40540 2858
rect 40788 800 40816 3538
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41052 3052 41104 3058
rect 41052 2994 41104 3000
rect 41064 800 41092 2994
rect 41340 800 41368 3470
rect 41880 2984 41932 2990
rect 41880 2926 41932 2932
rect 41604 2372 41656 2378
rect 41604 2314 41656 2320
rect 41616 800 41644 2314
rect 41892 800 41920 2926
rect 42168 800 42196 3606
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 42432 2508 42484 2514
rect 42432 2450 42484 2456
rect 42444 800 42472 2450
rect 42720 800 42748 3470
rect 42984 2916 43036 2922
rect 42984 2858 43036 2864
rect 42996 800 43024 2858
rect 43272 800 43300 3606
rect 44088 3596 44140 3602
rect 44088 3538 44140 3544
rect 43628 2848 43680 2854
rect 43548 2808 43628 2836
rect 43548 800 43576 2808
rect 43628 2790 43680 2796
rect 43812 2576 43864 2582
rect 43812 2518 43864 2524
rect 43824 800 43852 2518
rect 44100 800 44128 3538
rect 44916 3528 44968 3534
rect 44916 3470 44968 3476
rect 44364 2984 44416 2990
rect 44364 2926 44416 2932
rect 44376 800 44404 2926
rect 44640 2508 44692 2514
rect 44640 2450 44692 2456
rect 44652 800 44680 2450
rect 44928 800 44956 3470
rect 45192 2916 45244 2922
rect 45192 2858 45244 2864
rect 45204 800 45232 2858
rect 45480 800 45508 3606
rect 46296 3528 46348 3534
rect 46296 3470 46348 3476
rect 47124 3528 47176 3534
rect 47124 3470 47176 3476
rect 47676 3528 47728 3534
rect 47676 3470 47728 3476
rect 49056 3528 49108 3534
rect 49056 3470 49108 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 51540 3528 51592 3534
rect 51540 3470 51592 3476
rect 45744 2848 45796 2854
rect 45744 2790 45796 2796
rect 45756 800 45784 2790
rect 46020 2440 46072 2446
rect 46020 2382 46072 2388
rect 46032 800 46060 2382
rect 46308 800 46336 3470
rect 46572 2984 46624 2990
rect 46572 2926 46624 2932
rect 46584 800 46612 2926
rect 46848 2576 46900 2582
rect 46848 2518 46900 2524
rect 46860 800 46888 2518
rect 47136 800 47164 3470
rect 47400 2916 47452 2922
rect 47400 2858 47452 2864
rect 47412 800 47440 2858
rect 47688 800 47716 3470
rect 48780 2916 48832 2922
rect 48780 2858 48832 2864
rect 47952 2848 48004 2854
rect 47952 2790 48004 2796
rect 47964 800 47992 2790
rect 48228 2508 48280 2514
rect 48228 2450 48280 2456
rect 48240 800 48268 2450
rect 48504 2440 48556 2446
rect 48504 2382 48556 2388
rect 48516 800 48544 2382
rect 48792 800 48820 2858
rect 49068 800 49096 3470
rect 49332 2848 49384 2854
rect 49332 2790 49384 2796
rect 49344 800 49372 2790
rect 49620 800 49648 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 49884 2984 49936 2990
rect 49884 2926 49936 2932
rect 49896 800 49924 2926
rect 50712 2916 50764 2922
rect 50712 2858 50764 2864
rect 50160 2508 50212 2514
rect 50160 2450 50212 2456
rect 50172 800 50200 2450
rect 50620 2440 50672 2446
rect 50620 2382 50672 2388
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50632 1306 50660 2382
rect 50448 1278 50660 1306
rect 50448 800 50476 1278
rect 50724 800 50752 2858
rect 51000 800 51028 3470
rect 51264 2848 51316 2854
rect 51264 2790 51316 2796
rect 51276 800 51304 2790
rect 51552 800 51580 3470
rect 52092 2984 52144 2990
rect 52092 2926 52144 2932
rect 51816 2576 51868 2582
rect 51816 2518 51868 2524
rect 51828 800 51856 2518
rect 52104 800 52132 2926
rect 52368 2508 52420 2514
rect 52368 2450 52420 2456
rect 52380 800 52408 2450
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
<< via2 >>
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 12346 57452 12402 57488
rect 12346 57432 12348 57452
rect 12348 57432 12400 57452
rect 12400 57432 12402 57452
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 25686 56208 25742 56264
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 26330 56788 26332 56808
rect 26332 56788 26384 56808
rect 26384 56788 26386 56808
rect 26330 56752 26386 56788
rect 26514 56752 26570 56808
rect 27710 57432 27766 57488
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 29274 56344 29330 56400
rect 29826 57044 29882 57080
rect 29826 57024 29828 57044
rect 29828 57024 29880 57044
rect 29880 57024 29882 57044
rect 29550 56652 29552 56672
rect 29552 56652 29604 56672
rect 29604 56652 29606 56672
rect 29550 56616 29606 56652
rect 29826 56072 29882 56128
rect 32310 56788 32312 56808
rect 32312 56788 32364 56808
rect 32364 56788 32366 56808
rect 32310 56752 32366 56788
rect 32218 56072 32274 56128
rect 32678 55256 32734 55312
rect 33690 56788 33692 56808
rect 33692 56788 33744 56808
rect 33744 56788 33746 56808
rect 33690 56752 33746 56788
rect 34518 56652 34520 56672
rect 34520 56652 34572 56672
rect 34572 56652 34574 56672
rect 34518 56616 34574 56652
rect 34702 57044 34758 57080
rect 34702 57024 34704 57044
rect 34704 57024 34756 57044
rect 34756 57024 34758 57044
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 36082 56344 36138 56400
rect 35990 55256 36046 55312
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 37554 55936 37610 55992
rect 38382 55936 38438 55992
rect 39118 56480 39174 56536
rect 40774 56788 40776 56808
rect 40776 56788 40828 56808
rect 40828 56788 40830 56808
rect 40774 56752 40830 56788
rect 40590 56344 40646 56400
rect 41142 56924 41144 56944
rect 41144 56924 41196 56944
rect 41196 56924 41198 56944
rect 41142 56888 41198 56924
rect 41050 56072 41106 56128
rect 42246 56888 42302 56944
rect 41970 56788 41972 56808
rect 41972 56788 42024 56808
rect 42024 56788 42026 56808
rect 41970 56752 42026 56788
rect 41878 56228 41934 56264
rect 41878 56208 41880 56228
rect 41880 56208 41932 56228
rect 41932 56208 41934 56228
rect 44086 56788 44088 56808
rect 44088 56788 44140 56808
rect 44140 56788 44142 56808
rect 44086 56752 44142 56788
rect 44086 56208 44142 56264
rect 44270 55956 44326 55992
rect 44270 55936 44272 55956
rect 44272 55936 44324 55956
rect 44324 55936 44326 55956
rect 44822 56480 44878 56536
rect 45190 56344 45246 56400
rect 45834 56072 45890 56128
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 48686 56208 48742 56264
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
<< metal3 >>
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 12341 57490 12407 57493
rect 27705 57490 27771 57493
rect 12341 57488 27771 57490
rect 12341 57432 12346 57488
rect 12402 57432 27710 57488
rect 27766 57432 27771 57488
rect 12341 57430 27771 57432
rect 12341 57427 12407 57430
rect 27705 57427 27771 57430
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 29821 57082 29887 57085
rect 34697 57082 34763 57085
rect 29821 57080 34763 57082
rect 29821 57024 29826 57080
rect 29882 57024 34702 57080
rect 34758 57024 34763 57080
rect 29821 57022 34763 57024
rect 29821 57019 29887 57022
rect 34697 57019 34763 57022
rect 41137 56946 41203 56949
rect 42241 56946 42307 56949
rect 41137 56944 42307 56946
rect 41137 56888 41142 56944
rect 41198 56888 42246 56944
rect 42302 56888 42307 56944
rect 41137 56886 42307 56888
rect 41137 56883 41203 56886
rect 42241 56883 42307 56886
rect 26325 56810 26391 56813
rect 26509 56810 26575 56813
rect 26325 56808 26575 56810
rect 26325 56752 26330 56808
rect 26386 56752 26514 56808
rect 26570 56752 26575 56808
rect 26325 56750 26575 56752
rect 26325 56747 26391 56750
rect 26509 56747 26575 56750
rect 32305 56810 32371 56813
rect 33685 56810 33751 56813
rect 32305 56808 33751 56810
rect 32305 56752 32310 56808
rect 32366 56752 33690 56808
rect 33746 56752 33751 56808
rect 32305 56750 33751 56752
rect 32305 56747 32371 56750
rect 33685 56747 33751 56750
rect 40769 56810 40835 56813
rect 41965 56810 42031 56813
rect 44081 56810 44147 56813
rect 40769 56808 44147 56810
rect 40769 56752 40774 56808
rect 40830 56752 41970 56808
rect 42026 56752 44086 56808
rect 44142 56752 44147 56808
rect 40769 56750 44147 56752
rect 40769 56747 40835 56750
rect 41965 56747 42031 56750
rect 44081 56747 44147 56750
rect 29545 56674 29611 56677
rect 34513 56674 34579 56677
rect 29545 56672 34579 56674
rect 29545 56616 29550 56672
rect 29606 56616 34518 56672
rect 34574 56616 34579 56672
rect 29545 56614 34579 56616
rect 29545 56611 29611 56614
rect 34513 56611 34579 56614
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 39113 56538 39179 56541
rect 44817 56538 44883 56541
rect 39113 56536 44883 56538
rect 39113 56480 39118 56536
rect 39174 56480 44822 56536
rect 44878 56480 44883 56536
rect 39113 56478 44883 56480
rect 39113 56475 39179 56478
rect 44817 56475 44883 56478
rect 29269 56402 29335 56405
rect 36077 56402 36143 56405
rect 29269 56400 36143 56402
rect 29269 56344 29274 56400
rect 29330 56344 36082 56400
rect 36138 56344 36143 56400
rect 29269 56342 36143 56344
rect 29269 56339 29335 56342
rect 36077 56339 36143 56342
rect 40585 56402 40651 56405
rect 45185 56402 45251 56405
rect 40585 56400 45251 56402
rect 40585 56344 40590 56400
rect 40646 56344 45190 56400
rect 45246 56344 45251 56400
rect 40585 56342 45251 56344
rect 40585 56339 40651 56342
rect 45185 56339 45251 56342
rect 25681 56266 25747 56269
rect 41873 56266 41939 56269
rect 25681 56264 41939 56266
rect 25681 56208 25686 56264
rect 25742 56208 41878 56264
rect 41934 56208 41939 56264
rect 25681 56206 41939 56208
rect 25681 56203 25747 56206
rect 41873 56203 41939 56206
rect 44081 56266 44147 56269
rect 48681 56266 48747 56269
rect 44081 56264 48747 56266
rect 44081 56208 44086 56264
rect 44142 56208 48686 56264
rect 48742 56208 48747 56264
rect 44081 56206 48747 56208
rect 44081 56203 44147 56206
rect 48681 56203 48747 56206
rect 29821 56130 29887 56133
rect 32213 56130 32279 56133
rect 29821 56128 32279 56130
rect 29821 56072 29826 56128
rect 29882 56072 32218 56128
rect 32274 56072 32279 56128
rect 29821 56070 32279 56072
rect 29821 56067 29887 56070
rect 32213 56067 32279 56070
rect 41045 56130 41111 56133
rect 45829 56130 45895 56133
rect 41045 56128 45895 56130
rect 41045 56072 41050 56128
rect 41106 56072 45834 56128
rect 45890 56072 45895 56128
rect 41045 56070 45895 56072
rect 41045 56067 41111 56070
rect 45829 56067 45895 56070
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 37549 55994 37615 55997
rect 38377 55994 38443 55997
rect 44265 55994 44331 55997
rect 37549 55992 44331 55994
rect 37549 55936 37554 55992
rect 37610 55936 38382 55992
rect 38438 55936 44270 55992
rect 44326 55936 44331 55992
rect 37549 55934 44331 55936
rect 37549 55931 37615 55934
rect 38377 55931 38443 55934
rect 44265 55931 44331 55934
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 32673 55314 32739 55317
rect 35985 55314 36051 55317
rect 32673 55312 36051 55314
rect 32673 55256 32678 55312
rect 32734 55256 35990 55312
rect 36046 55256 36051 55312
rect 32673 55254 36051 55256
rect 32673 55251 32739 55254
rect 35985 55251 36051 55254
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23092 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1666464484
transform -1 0 26036 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1666464484
transform -1 0 32568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1666464484
transform 1 0 30268 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1666464484
transform 1 0 26312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1666464484
transform 1 0 26404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A_N
timestamp 1666464484
transform -1 0 35144 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B
timestamp 1666464484
transform 1 0 36248 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__B1
timestamp 1666464484
transform -1 0 29440 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A_N
timestamp 1666464484
transform 1 0 46092 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__B1
timestamp 1666464484
transform -1 0 38640 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B1
timestamp 1666464484
transform -1 0 27416 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1666464484
transform 1 0 35696 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__B2
timestamp 1666464484
transform 1 0 37260 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A2
timestamp 1666464484
transform 1 0 34868 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1666464484
transform 1 0 40204 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A2
timestamp 1666464484
transform -1 0 41124 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1666464484
transform 1 0 23920 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1666464484
transform 1 0 24472 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A2
timestamp 1666464484
transform 1 0 37628 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A2
timestamp 1666464484
transform 1 0 39376 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A1
timestamp 1666464484
transform 1 0 33580 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A1
timestamp 1666464484
transform 1 0 42688 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1666464484
transform -1 0 23552 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1666464484
transform 1 0 24472 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A1
timestamp 1666464484
transform 1 0 33580 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1666464484
transform 1 0 30360 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B1
timestamp 1666464484
transform 1 0 31280 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A1
timestamp 1666464484
transform 1 0 31832 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__B1
timestamp 1666464484
transform -1 0 40020 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A1
timestamp 1666464484
transform 1 0 41308 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A
timestamp 1666464484
transform -1 0 26588 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1666464484
transform 1 0 26404 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1666464484
transform -1 0 28888 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A2
timestamp 1666464484
transform -1 0 33212 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A2
timestamp 1666464484
transform 1 0 37260 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A1
timestamp 1666464484
transform 1 0 30176 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__C1
timestamp 1666464484
transform 1 0 28152 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 3772 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 27968 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 33304 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 37628 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 36984 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 42136 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 36156 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 42412 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666464484
transform -1 0 39192 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666464484
transform -1 0 40940 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666464484
transform -1 0 47012 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1666464484
transform -1 0 43700 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1666464484
transform -1 0 45724 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1666464484
transform -1 0 49220 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1666464484
transform -1 0 47748 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1666464484
transform -1 0 48392 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1666464484
transform -1 0 50324 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1666464484
transform -1 0 51612 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1666464484
transform -1 0 52992 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1666464484
transform -1 0 53912 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1666464484
transform -1 0 55660 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output22_A
timestamp 1666464484
transform 1 0 7176 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1666464484
transform 1 0 12236 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22
timestamp 1666464484
transform 1 0 3128 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4232 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43
timestamp 1666464484
transform 1 0 5060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55
timestamp 1666464484
transform 1 0 6164 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64
timestamp 1666464484
transform 1 0 6992 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1666464484
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1666464484
transform 1 0 10580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106
timestamp 1666464484
transform 1 0 10856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1666464484
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_124
timestamp 1666464484
transform 1 0 12512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_127
timestamp 1666464484
transform 1 0 12788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_138
timestamp 1666464484
transform 1 0 13800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1666464484
transform 1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_148
timestamp 1666464484
transform 1 0 14720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_159
timestamp 1666464484
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1666464484
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_180
timestamp 1666464484
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1666464484
transform 1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_190
timestamp 1666464484
transform 1 0 18584 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_201
timestamp 1666464484
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_208
timestamp 1666464484
transform 1 0 20240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_211
timestamp 1666464484
transform 1 0 20516 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_222
timestamp 1666464484
transform 1 0 21528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_229
timestamp 1666464484
transform 1 0 22172 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_232
timestamp 1666464484
transform 1 0 22448 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1666464484
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1666464484
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_264
timestamp 1666464484
transform 1 0 25392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1666464484
transform 1 0 26036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_274
timestamp 1666464484
transform 1 0 26312 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_285
timestamp 1666464484
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_292
timestamp 1666464484
transform 1 0 27968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_295
timestamp 1666464484
transform 1 0 28244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_306
timestamp 1666464484
transform 1 0 29256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_313
timestamp 1666464484
transform 1 0 29900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_316
timestamp 1666464484
transform 1 0 30176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1666464484
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1666464484
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_342
timestamp 1666464484
transform 1 0 32568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_349
timestamp 1666464484
transform 1 0 33212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_358
timestamp 1666464484
transform 1 0 34040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_363
timestamp 1666464484
transform 1 0 34500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_370
timestamp 1666464484
transform 1 0 35144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_379
timestamp 1666464484
transform 1 0 35972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_384
timestamp 1666464484
transform 1 0 36432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_391
timestamp 1666464484
transform 1 0 37076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_400
timestamp 1666464484
transform 1 0 37904 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_405
timestamp 1666464484
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1666464484
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1666464484
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_426
timestamp 1666464484
transform 1 0 40296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_433
timestamp 1666464484
transform 1 0 40940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_442
timestamp 1666464484
transform 1 0 41768 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_447
timestamp 1666464484
transform 1 0 42228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_454
timestamp 1666464484
transform 1 0 42872 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_463
timestamp 1666464484
transform 1 0 43700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_468
timestamp 1666464484
transform 1 0 44160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_475
timestamp 1666464484
transform 1 0 44804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_484
timestamp 1666464484
transform 1 0 45632 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1666464484
transform 1 0 46092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_496
timestamp 1666464484
transform 1 0 46736 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1666464484
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_510
timestamp 1666464484
transform 1 0 48024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_517
timestamp 1666464484
transform 1 0 48668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_526
timestamp 1666464484
transform 1 0 49496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_531
timestamp 1666464484
transform 1 0 49956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_538
timestamp 1666464484
transform 1 0 50600 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_547
timestamp 1666464484
transform 1 0 51428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_552
timestamp 1666464484
transform 1 0 51888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_559
timestamp 1666464484
transform 1 0 52532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_568
timestamp 1666464484
transform 1 0 53360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_573
timestamp 1666464484
transform 1 0 53820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_580
timestamp 1666464484
transform 1 0 54464 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1666464484
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_601
timestamp 1666464484
transform 1 0 56396 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_610
timestamp 1666464484
transform 1 0 57224 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_622 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 58328 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_44
timestamp 1666464484
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_56
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_64
timestamp 1666464484
transform 1 0 6992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_70
timestamp 1666464484
transform 1 0 7544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_77
timestamp 1666464484
transform 1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_84
timestamp 1666464484
transform 1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_87
timestamp 1666464484
transform 1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_92
timestamp 1666464484
transform 1 0 9568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_99
timestamp 1666464484
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_106
timestamp 1666464484
transform 1 0 10856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_120
timestamp 1666464484
transform 1 0 12144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_127
timestamp 1666464484
transform 1 0 12788 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_130
timestamp 1666464484
transform 1 0 13064 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_135
timestamp 1666464484
transform 1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1666464484
transform 1 0 14168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1666464484
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1666464484
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_170
timestamp 1666464484
transform 1 0 16744 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_173
timestamp 1666464484
transform 1 0 17020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1666464484
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_185
timestamp 1666464484
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1666464484
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_199
timestamp 1666464484
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_206
timestamp 1666464484
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_213
timestamp 1666464484
transform 1 0 20700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_216
timestamp 1666464484
transform 1 0 20976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_220 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21344 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_224
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_231
timestamp 1666464484
transform 1 0 22356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_256
timestamp 1666464484
transform 1 0 24656 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_259
timestamp 1666464484
transform 1 0 24932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_263
timestamp 1666464484
transform 1 0 25300 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_267
timestamp 1666464484
transform 1 0 25668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_274
timestamp 1666464484
transform 1 0 26312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_299
timestamp 1666464484
transform 1 0 28612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_302
timestamp 1666464484
transform 1 0 28888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_306
timestamp 1666464484
transform 1 0 29256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_310
timestamp 1666464484
transform 1 0 29624 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_314
timestamp 1666464484
transform 1 0 29992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_336
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_345
timestamp 1666464484
transform 1 0 32844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_368
timestamp 1666464484
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_375
timestamp 1666464484
transform 1 0 35604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_382
timestamp 1666464484
transform 1 0 36248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_386
timestamp 1666464484
transform 1 0 36616 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_388
timestamp 1666464484
transform 1 0 36800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_411
timestamp 1666464484
transform 1 0 38916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_418
timestamp 1666464484
transform 1 0 39560 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_425
timestamp 1666464484
transform 1 0 40204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_429
timestamp 1666464484
transform 1 0 40572 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_431
timestamp 1666464484
transform 1 0 40756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_436
timestamp 1666464484
transform 1 0 41216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_443
timestamp 1666464484
transform 1 0 41860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_450
timestamp 1666464484
transform 1 0 42504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_457
timestamp 1666464484
transform 1 0 43148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_464
timestamp 1666464484
transform 1 0 43792 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_471
timestamp 1666464484
transform 1 0 44436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_474
timestamp 1666464484
transform 1 0 44712 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_479
timestamp 1666464484
transform 1 0 45172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_486
timestamp 1666464484
transform 1 0 45816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_493
timestamp 1666464484
transform 1 0 46460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1666464484
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_507
timestamp 1666464484
transform 1 0 47748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_514
timestamp 1666464484
transform 1 0 48392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_517
timestamp 1666464484
transform 1 0 48668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_522
timestamp 1666464484
transform 1 0 49128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_529
timestamp 1666464484
transform 1 0 49772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_536
timestamp 1666464484
transform 1 0 50416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_543
timestamp 1666464484
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_550
timestamp 1666464484
transform 1 0 51704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_557
timestamp 1666464484
transform 1 0 52348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_560
timestamp 1666464484
transform 1 0 52624 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_565
timestamp 1666464484
transform 1 0 53084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_577
timestamp 1666464484
transform 1 0 54188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_589
timestamp 1666464484
transform 1 0 55292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_601
timestamp 1666464484
transform 1 0 56396 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_603
timestamp 1666464484
transform 1 0 56580 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_615
timestamp 1666464484
transform 1 0 57684 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_623
timestamp 1666464484
transform 1 0 58420 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_22
timestamp 1666464484
transform 1 0 3128 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_34
timestamp 1666464484
transform 1 0 4232 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_46
timestamp 1666464484
transform 1 0 5336 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_58
timestamp 1666464484
transform 1 0 6440 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1666464484
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_93
timestamp 1666464484
transform 1 0 9660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_99
timestamp 1666464484
transform 1 0 10212 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_103
timestamp 1666464484
transform 1 0 10580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_108
timestamp 1666464484
transform 1 0 11040 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1666464484
transform 1 0 11776 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_130
timestamp 1666464484
transform 1 0 13064 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_148
timestamp 1666464484
transform 1 0 14720 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1666464484
transform 1 0 14996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_156
timestamp 1666464484
transform 1 0 15456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 1666464484
transform 1 0 16100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_170
timestamp 1666464484
transform 1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1666464484
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_191
timestamp 1666464484
transform 1 0 18676 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_194
timestamp 1666464484
transform 1 0 18952 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_198
timestamp 1666464484
transform 1 0 19320 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1666464484
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_234
timestamp 1666464484
transform 1 0 22632 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_237
timestamp 1666464484
transform 1 0 22908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_241
timestamp 1666464484
transform 1 0 23276 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_245
timestamp 1666464484
transform 1 0 23644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_252
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_277
timestamp 1666464484
transform 1 0 26588 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_280
timestamp 1666464484
transform 1 0 26864 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_284
timestamp 1666464484
transform 1 0 27232 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_288
timestamp 1666464484
transform 1 0 27600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1666464484
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_320
timestamp 1666464484
transform 1 0 30544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_323
timestamp 1666464484
transform 1 0 30820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_328
timestamp 1666464484
transform 1 0 31280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_355
timestamp 1666464484
transform 1 0 33764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_362
timestamp 1666464484
transform 1 0 34408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_366
timestamp 1666464484
transform 1 0 34776 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_389
timestamp 1666464484
transform 1 0 36892 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_396
timestamp 1666464484
transform 1 0 37536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1666464484
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_407
timestamp 1666464484
transform 1 0 38548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_409
timestamp 1666464484
transform 1 0 38732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_414
timestamp 1666464484
transform 1 0 39192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_421
timestamp 1666464484
transform 1 0 39836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_428
timestamp 1666464484
transform 1 0 40480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_435
timestamp 1666464484
transform 1 0 41124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_442
timestamp 1666464484
transform 1 0 41768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_449
timestamp 1666464484
transform 1 0 42412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_452
timestamp 1666464484
transform 1 0 42688 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_457
timestamp 1666464484
transform 1 0 43148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_464
timestamp 1666464484
transform 1 0 43792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_471
timestamp 1666464484
transform 1 0 44436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_478
timestamp 1666464484
transform 1 0 45080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_485
timestamp 1666464484
transform 1 0 45724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_492
timestamp 1666464484
transform 1 0 46368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_495
timestamp 1666464484
transform 1 0 46644 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_500
timestamp 1666464484
transform 1 0 47104 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_507
timestamp 1666464484
transform 1 0 47748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_514
timestamp 1666464484
transform 1 0 48392 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_525
timestamp 1666464484
transform 1 0 49404 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_532
timestamp 1666464484
transform 1 0 50048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_536
timestamp 1666464484
transform 1 0 50416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_538
timestamp 1666464484
transform 1 0 50600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_542
timestamp 1666464484
transform 1 0 50968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_546
timestamp 1666464484
transform 1 0 51336 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_553
timestamp 1666464484
transform 1 0 51980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_565
timestamp 1666464484
transform 1 0 53084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_577
timestamp 1666464484
transform 1 0 54188 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_581
timestamp 1666464484
transform 1 0 54556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_593
timestamp 1666464484
transform 1 0 55660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_605
timestamp 1666464484
transform 1 0 56764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_617
timestamp 1666464484
transform 1 0 57868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_624
timestamp 1666464484
transform 1 0 58512 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_39
timestamp 1666464484
transform 1 0 4692 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1666464484
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_56
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_68
timestamp 1666464484
transform 1 0 7360 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_80
timestamp 1666464484
transform 1 0 8464 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_87
timestamp 1666464484
transform 1 0 9108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_99
timestamp 1666464484
transform 1 0 10212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_123
timestamp 1666464484
transform 1 0 12420 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_130
timestamp 1666464484
transform 1 0 13064 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_142
timestamp 1666464484
transform 1 0 14168 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_154
timestamp 1666464484
transform 1 0 15272 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_173
timestamp 1666464484
transform 1 0 17020 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_179
timestamp 1666464484
transform 1 0 17572 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_183
timestamp 1666464484
transform 1 0 17940 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_192
timestamp 1666464484
transform 1 0 18768 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_199
timestamp 1666464484
transform 1 0 19412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_206
timestamp 1666464484
transform 1 0 20056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_213
timestamp 1666464484
transform 1 0 20700 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_216
timestamp 1666464484
transform 1 0 20976 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_220
timestamp 1666464484
transform 1 0 21344 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_224
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_231
timestamp 1666464484
transform 1 0 22356 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_256
timestamp 1666464484
transform 1 0 24656 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_259
timestamp 1666464484
transform 1 0 24932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_263
timestamp 1666464484
transform 1 0 25300 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_267
timestamp 1666464484
transform 1 0 25668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_274
timestamp 1666464484
transform 1 0 26312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_299
timestamp 1666464484
transform 1 0 28612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_302
timestamp 1666464484
transform 1 0 28888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_306
timestamp 1666464484
transform 1 0 29256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_310
timestamp 1666464484
transform 1 0 29624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_317
timestamp 1666464484
transform 1 0 30268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_342
timestamp 1666464484
transform 1 0 32568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_345
timestamp 1666464484
transform 1 0 32844 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_368
timestamp 1666464484
transform 1 0 34960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_375
timestamp 1666464484
transform 1 0 35604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_382
timestamp 1666464484
transform 1 0 36248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_386
timestamp 1666464484
transform 1 0 36616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_388
timestamp 1666464484
transform 1 0 36800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_411
timestamp 1666464484
transform 1 0 38916 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_418
timestamp 1666464484
transform 1 0 39560 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_425
timestamp 1666464484
transform 1 0 40204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_429
timestamp 1666464484
transform 1 0 40572 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_431
timestamp 1666464484
transform 1 0 40756 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_436
timestamp 1666464484
transform 1 0 41216 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_448
timestamp 1666464484
transform 1 0 42320 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_460
timestamp 1666464484
transform 1 0 43424 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_472
timestamp 1666464484
transform 1 0 44528 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_474
timestamp 1666464484
transform 1 0 44712 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_486
timestamp 1666464484
transform 1 0 45816 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_498
timestamp 1666464484
transform 1 0 46920 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_510
timestamp 1666464484
transform 1 0 48024 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1666464484
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1666464484
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1666464484
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1666464484
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_560
timestamp 1666464484
transform 1 0 52624 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_572
timestamp 1666464484
transform 1 0 53728 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_584
timestamp 1666464484
transform 1 0 54832 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_596
timestamp 1666464484
transform 1 0 55936 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_603
timestamp 1666464484
transform 1 0 56580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_615
timestamp 1666464484
transform 1 0 57684 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_623
timestamp 1666464484
transform 1 0 58420 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_22
timestamp 1666464484
transform 1 0 3128 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_34
timestamp 1666464484
transform 1 0 4232 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_46
timestamp 1666464484
transform 1 0 5336 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_58
timestamp 1666464484
transform 1 0 6440 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_89
timestamp 1666464484
transform 1 0 9292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_101
timestamp 1666464484
transform 1 0 10396 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_108
timestamp 1666464484
transform 1 0 11040 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_120
timestamp 1666464484
transform 1 0 12144 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_132
timestamp 1666464484
transform 1 0 13248 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_144
timestamp 1666464484
transform 1 0 14352 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_151
timestamp 1666464484
transform 1 0 14996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_163
timestamp 1666464484
transform 1 0 16100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_175
timestamp 1666464484
transform 1 0 17204 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_187
timestamp 1666464484
transform 1 0 18308 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_194
timestamp 1666464484
transform 1 0 18952 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_201
timestamp 1666464484
transform 1 0 19596 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_213
timestamp 1666464484
transform 1 0 20700 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_220
timestamp 1666464484
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_227
timestamp 1666464484
transform 1 0 21988 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_234
timestamp 1666464484
transform 1 0 22632 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_237
timestamp 1666464484
transform 1 0 22908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_241
timestamp 1666464484
transform 1 0 23276 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_245
timestamp 1666464484
transform 1 0 23644 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_252
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_277
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_280
timestamp 1666464484
transform 1 0 26864 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_284
timestamp 1666464484
transform 1 0 27232 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_288
timestamp 1666464484
transform 1 0 27600 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_295
timestamp 1666464484
transform 1 0 28244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_320
timestamp 1666464484
transform 1 0 30544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_323
timestamp 1666464484
transform 1 0 30820 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_331
timestamp 1666464484
transform 1 0 31556 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_335
timestamp 1666464484
transform 1 0 31924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_357
timestamp 1666464484
transform 1 0 33948 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_366
timestamp 1666464484
transform 1 0 34776 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_389
timestamp 1666464484
transform 1 0 36892 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_396
timestamp 1666464484
transform 1 0 37536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1666464484
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_407
timestamp 1666464484
transform 1 0 38548 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_409
timestamp 1666464484
transform 1 0 38732 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_414
timestamp 1666464484
transform 1 0 39192 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_426
timestamp 1666464484
transform 1 0 40296 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_438
timestamp 1666464484
transform 1 0 41400 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_450
timestamp 1666464484
transform 1 0 42504 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_452
timestamp 1666464484
transform 1 0 42688 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_464
timestamp 1666464484
transform 1 0 43792 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_476
timestamp 1666464484
transform 1 0 44896 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_488
timestamp 1666464484
transform 1 0 46000 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_495
timestamp 1666464484
transform 1 0 46644 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_507
timestamp 1666464484
transform 1 0 47748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_519
timestamp 1666464484
transform 1 0 48852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_531
timestamp 1666464484
transform 1 0 49956 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_538
timestamp 1666464484
transform 1 0 50600 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_550
timestamp 1666464484
transform 1 0 51704 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_562
timestamp 1666464484
transform 1 0 52808 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_574
timestamp 1666464484
transform 1 0 53912 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_581
timestamp 1666464484
transform 1 0 54556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_593
timestamp 1666464484
transform 1 0 55660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_605
timestamp 1666464484
transform 1 0 56764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_617
timestamp 1666464484
transform 1 0 57868 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_624
timestamp 1666464484
transform 1 0 58512 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_39
timestamp 1666464484
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_44
timestamp 1666464484
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_56
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_68
timestamp 1666464484
transform 1 0 7360 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_80
timestamp 1666464484
transform 1 0 8464 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_87
timestamp 1666464484
transform 1 0 9108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_99
timestamp 1666464484
transform 1 0 10212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_123
timestamp 1666464484
transform 1 0 12420 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_130
timestamp 1666464484
transform 1 0 13064 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_142
timestamp 1666464484
transform 1 0 14168 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_154
timestamp 1666464484
transform 1 0 15272 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_166
timestamp 1666464484
transform 1 0 16376 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_173
timestamp 1666464484
transform 1 0 17020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_185
timestamp 1666464484
transform 1 0 18124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_197
timestamp 1666464484
transform 1 0 19228 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_209
timestamp 1666464484
transform 1 0 20332 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_216
timestamp 1666464484
transform 1 0 20976 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_231
timestamp 1666464484
transform 1 0 22356 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_256
timestamp 1666464484
transform 1 0 24656 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_259
timestamp 1666464484
transform 1 0 24932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_264
timestamp 1666464484
transform 1 0 25392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_274
timestamp 1666464484
transform 1 0 26312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_299
timestamp 1666464484
transform 1 0 28612 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_302
timestamp 1666464484
transform 1 0 28888 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_311
timestamp 1666464484
transform 1 0 29716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_336
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_342
timestamp 1666464484
transform 1 0 32568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_345
timestamp 1666464484
transform 1 0 32844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_369
timestamp 1666464484
transform 1 0 35052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_376
timestamp 1666464484
transform 1 0 35696 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_383
timestamp 1666464484
transform 1 0 36340 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_388
timestamp 1666464484
transform 1 0 36800 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_400
timestamp 1666464484
transform 1 0 37904 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_412
timestamp 1666464484
transform 1 0 39008 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_424
timestamp 1666464484
transform 1 0 40112 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_431
timestamp 1666464484
transform 1 0 40756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_443
timestamp 1666464484
transform 1 0 41860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_455
timestamp 1666464484
transform 1 0 42964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_467
timestamp 1666464484
transform 1 0 44068 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_474
timestamp 1666464484
transform 1 0 44712 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_486
timestamp 1666464484
transform 1 0 45816 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_498
timestamp 1666464484
transform 1 0 46920 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_510
timestamp 1666464484
transform 1 0 48024 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1666464484
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1666464484
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1666464484
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1666464484
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_560
timestamp 1666464484
transform 1 0 52624 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_572
timestamp 1666464484
transform 1 0 53728 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_584
timestamp 1666464484
transform 1 0 54832 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_596
timestamp 1666464484
transform 1 0 55936 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_603
timestamp 1666464484
transform 1 0 56580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_615
timestamp 1666464484
transform 1 0 57684 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_623
timestamp 1666464484
transform 1 0 58420 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_22
timestamp 1666464484
transform 1 0 3128 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_34
timestamp 1666464484
transform 1 0 4232 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_46
timestamp 1666464484
transform 1 0 5336 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_58
timestamp 1666464484
transform 1 0 6440 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_89
timestamp 1666464484
transform 1 0 9292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_101
timestamp 1666464484
transform 1 0 10396 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_108
timestamp 1666464484
transform 1 0 11040 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_120
timestamp 1666464484
transform 1 0 12144 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_132
timestamp 1666464484
transform 1 0 13248 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_144
timestamp 1666464484
transform 1 0 14352 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_151
timestamp 1666464484
transform 1 0 14996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_163
timestamp 1666464484
transform 1 0 16100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_175
timestamp 1666464484
transform 1 0 17204 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_187
timestamp 1666464484
transform 1 0 18308 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_194
timestamp 1666464484
transform 1 0 18952 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_206
timestamp 1666464484
transform 1 0 20056 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_218
timestamp 1666464484
transform 1 0 21160 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_230
timestamp 1666464484
transform 1 0 22264 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_237
timestamp 1666464484
transform 1 0 22908 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_243
timestamp 1666464484
transform 1 0 23460 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_252
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_280
timestamp 1666464484
transform 1 0 26864 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_286
timestamp 1666464484
transform 1 0 27416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_308
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_320
timestamp 1666464484
transform 1 0 30544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_323
timestamp 1666464484
transform 1 0 30820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_346
timestamp 1666464484
transform 1 0 32936 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_353
timestamp 1666464484
transform 1 0 33580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1666464484
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_364
timestamp 1666464484
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_366
timestamp 1666464484
transform 1 0 34776 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_371
timestamp 1666464484
transform 1 0 35236 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_383
timestamp 1666464484
transform 1 0 36340 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_395
timestamp 1666464484
transform 1 0 37444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_407
timestamp 1666464484
transform 1 0 38548 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_409
timestamp 1666464484
transform 1 0 38732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1666464484
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1666464484
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_445
timestamp 1666464484
transform 1 0 42044 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_452
timestamp 1666464484
transform 1 0 42688 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_464
timestamp 1666464484
transform 1 0 43792 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_476
timestamp 1666464484
transform 1 0 44896 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_488
timestamp 1666464484
transform 1 0 46000 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_495
timestamp 1666464484
transform 1 0 46644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_507
timestamp 1666464484
transform 1 0 47748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_519
timestamp 1666464484
transform 1 0 48852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_531
timestamp 1666464484
transform 1 0 49956 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_538
timestamp 1666464484
transform 1 0 50600 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_550
timestamp 1666464484
transform 1 0 51704 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_562
timestamp 1666464484
transform 1 0 52808 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_574
timestamp 1666464484
transform 1 0 53912 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_581
timestamp 1666464484
transform 1 0 54556 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_593
timestamp 1666464484
transform 1 0 55660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_605
timestamp 1666464484
transform 1 0 56764 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_617
timestamp 1666464484
transform 1 0 57868 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_624
timestamp 1666464484
transform 1 0 58512 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_39
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_44
timestamp 1666464484
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_56
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_68
timestamp 1666464484
transform 1 0 7360 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_80
timestamp 1666464484
transform 1 0 8464 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_87
timestamp 1666464484
transform 1 0 9108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_99
timestamp 1666464484
transform 1 0 10212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_123
timestamp 1666464484
transform 1 0 12420 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_130
timestamp 1666464484
transform 1 0 13064 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_142
timestamp 1666464484
transform 1 0 14168 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_154
timestamp 1666464484
transform 1 0 15272 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_166
timestamp 1666464484
transform 1 0 16376 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_173
timestamp 1666464484
transform 1 0 17020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_185
timestamp 1666464484
transform 1 0 18124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_197
timestamp 1666464484
transform 1 0 19228 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_209
timestamp 1666464484
transform 1 0 20332 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_216
timestamp 1666464484
transform 1 0 20976 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_228
timestamp 1666464484
transform 1 0 22080 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_240
timestamp 1666464484
transform 1 0 23184 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_248
timestamp 1666464484
transform 1 0 23920 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_252
timestamp 1666464484
transform 1 0 24288 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_259
timestamp 1666464484
transform 1 0 24932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_263
timestamp 1666464484
transform 1 0 25300 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_267
timestamp 1666464484
transform 1 0 25668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_274
timestamp 1666464484
transform 1 0 26312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_299
timestamp 1666464484
transform 1 0 28612 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_302
timestamp 1666464484
transform 1 0 28888 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_308
timestamp 1666464484
transform 1 0 29440 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_330
timestamp 1666464484
transform 1 0 31464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_343
timestamp 1666464484
transform 1 0 32660 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_345
timestamp 1666464484
transform 1 0 32844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_350
timestamp 1666464484
transform 1 0 33304 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_356
timestamp 1666464484
transform 1 0 33856 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_378
timestamp 1666464484
transform 1 0 35880 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_386
timestamp 1666464484
transform 1 0 36616 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_388
timestamp 1666464484
transform 1 0 36800 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_400
timestamp 1666464484
transform 1 0 37904 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_412
timestamp 1666464484
transform 1 0 39008 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_424
timestamp 1666464484
transform 1 0 40112 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_431
timestamp 1666464484
transform 1 0 40756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_443
timestamp 1666464484
transform 1 0 41860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_455
timestamp 1666464484
transform 1 0 42964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_467
timestamp 1666464484
transform 1 0 44068 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_474
timestamp 1666464484
transform 1 0 44712 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_486
timestamp 1666464484
transform 1 0 45816 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_498
timestamp 1666464484
transform 1 0 46920 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_510
timestamp 1666464484
transform 1 0 48024 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1666464484
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1666464484
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1666464484
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1666464484
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_560
timestamp 1666464484
transform 1 0 52624 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_572
timestamp 1666464484
transform 1 0 53728 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_584
timestamp 1666464484
transform 1 0 54832 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_596
timestamp 1666464484
transform 1 0 55936 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_603
timestamp 1666464484
transform 1 0 56580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_615
timestamp 1666464484
transform 1 0 57684 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_623
timestamp 1666464484
transform 1 0 58420 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_22
timestamp 1666464484
transform 1 0 3128 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_34
timestamp 1666464484
transform 1 0 4232 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_46
timestamp 1666464484
transform 1 0 5336 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_58
timestamp 1666464484
transform 1 0 6440 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_89
timestamp 1666464484
transform 1 0 9292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_101
timestamp 1666464484
transform 1 0 10396 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_108
timestamp 1666464484
transform 1 0 11040 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_120
timestamp 1666464484
transform 1 0 12144 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_132
timestamp 1666464484
transform 1 0 13248 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_144
timestamp 1666464484
transform 1 0 14352 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_151
timestamp 1666464484
transform 1 0 14996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_163
timestamp 1666464484
transform 1 0 16100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_175
timestamp 1666464484
transform 1 0 17204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_187
timestamp 1666464484
transform 1 0 18308 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_194
timestamp 1666464484
transform 1 0 18952 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_206
timestamp 1666464484
transform 1 0 20056 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_218
timestamp 1666464484
transform 1 0 21160 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_230
timestamp 1666464484
transform 1 0 22264 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_237
timestamp 1666464484
transform 1 0 22908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_249
timestamp 1666464484
transform 1 0 24012 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_261
timestamp 1666464484
transform 1 0 25116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_267
timestamp 1666464484
transform 1 0 25668 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_271
timestamp 1666464484
transform 1 0 26036 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_277
timestamp 1666464484
transform 1 0 26588 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_280
timestamp 1666464484
transform 1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_284
timestamp 1666464484
transform 1 0 27232 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_288
timestamp 1666464484
transform 1 0 27600 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_313
timestamp 1666464484
transform 1 0 29900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_320
timestamp 1666464484
transform 1 0 30544 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_323
timestamp 1666464484
transform 1 0 30820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_328
timestamp 1666464484
transform 1 0 31280 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_336
timestamp 1666464484
transform 1 0 32016 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_340
timestamp 1666464484
transform 1 0 32384 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_352
timestamp 1666464484
transform 1 0 33488 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_364
timestamp 1666464484
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_366
timestamp 1666464484
transform 1 0 34776 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_378
timestamp 1666464484
transform 1 0 35880 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_390
timestamp 1666464484
transform 1 0 36984 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_402
timestamp 1666464484
transform 1 0 38088 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_409
timestamp 1666464484
transform 1 0 38732 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1666464484
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1666464484
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_445
timestamp 1666464484
transform 1 0 42044 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_452
timestamp 1666464484
transform 1 0 42688 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_464
timestamp 1666464484
transform 1 0 43792 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_476
timestamp 1666464484
transform 1 0 44896 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_488
timestamp 1666464484
transform 1 0 46000 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_495
timestamp 1666464484
transform 1 0 46644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_507
timestamp 1666464484
transform 1 0 47748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_519
timestamp 1666464484
transform 1 0 48852 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_531
timestamp 1666464484
transform 1 0 49956 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_538
timestamp 1666464484
transform 1 0 50600 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_550
timestamp 1666464484
transform 1 0 51704 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_562
timestamp 1666464484
transform 1 0 52808 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_574
timestamp 1666464484
transform 1 0 53912 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_581
timestamp 1666464484
transform 1 0 54556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_593
timestamp 1666464484
transform 1 0 55660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_605
timestamp 1666464484
transform 1 0 56764 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_617
timestamp 1666464484
transform 1 0 57868 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_624
timestamp 1666464484
transform 1 0 58512 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_39
timestamp 1666464484
transform 1 0 4692 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1666464484
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_56
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_68
timestamp 1666464484
transform 1 0 7360 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_80
timestamp 1666464484
transform 1 0 8464 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_87
timestamp 1666464484
transform 1 0 9108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_99
timestamp 1666464484
transform 1 0 10212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_123
timestamp 1666464484
transform 1 0 12420 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_130
timestamp 1666464484
transform 1 0 13064 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_142
timestamp 1666464484
transform 1 0 14168 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_154
timestamp 1666464484
transform 1 0 15272 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_166
timestamp 1666464484
transform 1 0 16376 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_173
timestamp 1666464484
transform 1 0 17020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_185
timestamp 1666464484
transform 1 0 18124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_197
timestamp 1666464484
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_209
timestamp 1666464484
transform 1 0 20332 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_216
timestamp 1666464484
transform 1 0 20976 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_228
timestamp 1666464484
transform 1 0 22080 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_240
timestamp 1666464484
transform 1 0 23184 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_252
timestamp 1666464484
transform 1 0 24288 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_259
timestamp 1666464484
transform 1 0 24932 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_267
timestamp 1666464484
transform 1 0 25668 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_289
timestamp 1666464484
transform 1 0 27692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_296
timestamp 1666464484
transform 1 0 28336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_300
timestamp 1666464484
transform 1 0 28704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_302
timestamp 1666464484
transform 1 0 28888 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_313
timestamp 1666464484
transform 1 0 29900 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_319
timestamp 1666464484
transform 1 0 30452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_331
timestamp 1666464484
transform 1 0 31556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_343
timestamp 1666464484
transform 1 0 32660 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_345
timestamp 1666464484
transform 1 0 32844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_357
timestamp 1666464484
transform 1 0 33948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_369
timestamp 1666464484
transform 1 0 35052 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_381
timestamp 1666464484
transform 1 0 36156 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_388
timestamp 1666464484
transform 1 0 36800 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_400
timestamp 1666464484
transform 1 0 37904 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_412
timestamp 1666464484
transform 1 0 39008 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_424
timestamp 1666464484
transform 1 0 40112 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_431
timestamp 1666464484
transform 1 0 40756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_443
timestamp 1666464484
transform 1 0 41860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_455
timestamp 1666464484
transform 1 0 42964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_467
timestamp 1666464484
transform 1 0 44068 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_474
timestamp 1666464484
transform 1 0 44712 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_486
timestamp 1666464484
transform 1 0 45816 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_498
timestamp 1666464484
transform 1 0 46920 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_510
timestamp 1666464484
transform 1 0 48024 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1666464484
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1666464484
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1666464484
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1666464484
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_560
timestamp 1666464484
transform 1 0 52624 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_572
timestamp 1666464484
transform 1 0 53728 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_584
timestamp 1666464484
transform 1 0 54832 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_596
timestamp 1666464484
transform 1 0 55936 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_603
timestamp 1666464484
transform 1 0 56580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_615
timestamp 1666464484
transform 1 0 57684 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_623
timestamp 1666464484
transform 1 0 58420 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_15
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_22
timestamp 1666464484
transform 1 0 3128 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_34
timestamp 1666464484
transform 1 0 4232 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_46
timestamp 1666464484
transform 1 0 5336 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_58
timestamp 1666464484
transform 1 0 6440 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_89
timestamp 1666464484
transform 1 0 9292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_101
timestamp 1666464484
transform 1 0 10396 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_108
timestamp 1666464484
transform 1 0 11040 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_120
timestamp 1666464484
transform 1 0 12144 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_132
timestamp 1666464484
transform 1 0 13248 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_144
timestamp 1666464484
transform 1 0 14352 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_151
timestamp 1666464484
transform 1 0 14996 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_163
timestamp 1666464484
transform 1 0 16100 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_175
timestamp 1666464484
transform 1 0 17204 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_187
timestamp 1666464484
transform 1 0 18308 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_194
timestamp 1666464484
transform 1 0 18952 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_206
timestamp 1666464484
transform 1 0 20056 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_218
timestamp 1666464484
transform 1 0 21160 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_230
timestamp 1666464484
transform 1 0 22264 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_237
timestamp 1666464484
transform 1 0 22908 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_249
timestamp 1666464484
transform 1 0 24012 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_261
timestamp 1666464484
transform 1 0 25116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_273
timestamp 1666464484
transform 1 0 26220 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_276
timestamp 1666464484
transform 1 0 26496 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_280
timestamp 1666464484
transform 1 0 26864 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_292
timestamp 1666464484
transform 1 0 27968 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_304
timestamp 1666464484
transform 1 0 29072 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_316
timestamp 1666464484
transform 1 0 30176 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_323
timestamp 1666464484
transform 1 0 30820 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_335
timestamp 1666464484
transform 1 0 31924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_347
timestamp 1666464484
transform 1 0 33028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_359
timestamp 1666464484
transform 1 0 34132 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_366
timestamp 1666464484
transform 1 0 34776 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_378
timestamp 1666464484
transform 1 0 35880 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_390
timestamp 1666464484
transform 1 0 36984 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_402
timestamp 1666464484
transform 1 0 38088 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_409
timestamp 1666464484
transform 1 0 38732 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1666464484
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1666464484
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_445
timestamp 1666464484
transform 1 0 42044 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_452
timestamp 1666464484
transform 1 0 42688 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_464
timestamp 1666464484
transform 1 0 43792 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_476
timestamp 1666464484
transform 1 0 44896 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_488
timestamp 1666464484
transform 1 0 46000 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_495
timestamp 1666464484
transform 1 0 46644 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_507
timestamp 1666464484
transform 1 0 47748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_519
timestamp 1666464484
transform 1 0 48852 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_531
timestamp 1666464484
transform 1 0 49956 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_538
timestamp 1666464484
transform 1 0 50600 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_550
timestamp 1666464484
transform 1 0 51704 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_562
timestamp 1666464484
transform 1 0 52808 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_574
timestamp 1666464484
transform 1 0 53912 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_581
timestamp 1666464484
transform 1 0 54556 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_593
timestamp 1666464484
transform 1 0 55660 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_605
timestamp 1666464484
transform 1 0 56764 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_617
timestamp 1666464484
transform 1 0 57868 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_624
timestamp 1666464484
transform 1 0 58512 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_44
timestamp 1666464484
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_56
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_68
timestamp 1666464484
transform 1 0 7360 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_80
timestamp 1666464484
transform 1 0 8464 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_87
timestamp 1666464484
transform 1 0 9108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_99
timestamp 1666464484
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_123
timestamp 1666464484
transform 1 0 12420 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_130
timestamp 1666464484
transform 1 0 13064 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_142
timestamp 1666464484
transform 1 0 14168 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_154
timestamp 1666464484
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_166
timestamp 1666464484
transform 1 0 16376 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_173
timestamp 1666464484
transform 1 0 17020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_185
timestamp 1666464484
transform 1 0 18124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_197
timestamp 1666464484
transform 1 0 19228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_209
timestamp 1666464484
transform 1 0 20332 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_216
timestamp 1666464484
transform 1 0 20976 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_228
timestamp 1666464484
transform 1 0 22080 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_240
timestamp 1666464484
transform 1 0 23184 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_252
timestamp 1666464484
transform 1 0 24288 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_259
timestamp 1666464484
transform 1 0 24932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_271
timestamp 1666464484
transform 1 0 26036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_283
timestamp 1666464484
transform 1 0 27140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_295
timestamp 1666464484
transform 1 0 28244 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_302
timestamp 1666464484
transform 1 0 28888 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_314
timestamp 1666464484
transform 1 0 29992 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_326
timestamp 1666464484
transform 1 0 31096 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_338
timestamp 1666464484
transform 1 0 32200 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_345
timestamp 1666464484
transform 1 0 32844 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_357
timestamp 1666464484
transform 1 0 33948 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_369
timestamp 1666464484
transform 1 0 35052 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_381
timestamp 1666464484
transform 1 0 36156 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_388
timestamp 1666464484
transform 1 0 36800 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_400
timestamp 1666464484
transform 1 0 37904 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_412
timestamp 1666464484
transform 1 0 39008 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_424
timestamp 1666464484
transform 1 0 40112 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_431
timestamp 1666464484
transform 1 0 40756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_443
timestamp 1666464484
transform 1 0 41860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_455
timestamp 1666464484
transform 1 0 42964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_467
timestamp 1666464484
transform 1 0 44068 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_474
timestamp 1666464484
transform 1 0 44712 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_486
timestamp 1666464484
transform 1 0 45816 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_498
timestamp 1666464484
transform 1 0 46920 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_510
timestamp 1666464484
transform 1 0 48024 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1666464484
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1666464484
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1666464484
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1666464484
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_560
timestamp 1666464484
transform 1 0 52624 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_572
timestamp 1666464484
transform 1 0 53728 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_584
timestamp 1666464484
transform 1 0 54832 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_596
timestamp 1666464484
transform 1 0 55936 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_603
timestamp 1666464484
transform 1 0 56580 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_615
timestamp 1666464484
transform 1 0 57684 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_623
timestamp 1666464484
transform 1 0 58420 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_22
timestamp 1666464484
transform 1 0 3128 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_34
timestamp 1666464484
transform 1 0 4232 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_46
timestamp 1666464484
transform 1 0 5336 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_58
timestamp 1666464484
transform 1 0 6440 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_89
timestamp 1666464484
transform 1 0 9292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_101
timestamp 1666464484
transform 1 0 10396 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_108
timestamp 1666464484
transform 1 0 11040 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_120
timestamp 1666464484
transform 1 0 12144 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_132
timestamp 1666464484
transform 1 0 13248 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_144
timestamp 1666464484
transform 1 0 14352 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_151
timestamp 1666464484
transform 1 0 14996 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_163
timestamp 1666464484
transform 1 0 16100 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_175
timestamp 1666464484
transform 1 0 17204 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_187
timestamp 1666464484
transform 1 0 18308 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_194
timestamp 1666464484
transform 1 0 18952 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_206
timestamp 1666464484
transform 1 0 20056 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_218
timestamp 1666464484
transform 1 0 21160 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_230
timestamp 1666464484
transform 1 0 22264 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_237
timestamp 1666464484
transform 1 0 22908 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_249
timestamp 1666464484
transform 1 0 24012 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_261
timestamp 1666464484
transform 1 0 25116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_273
timestamp 1666464484
transform 1 0 26220 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_280
timestamp 1666464484
transform 1 0 26864 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_292
timestamp 1666464484
transform 1 0 27968 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_304
timestamp 1666464484
transform 1 0 29072 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_316
timestamp 1666464484
transform 1 0 30176 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_323
timestamp 1666464484
transform 1 0 30820 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_335
timestamp 1666464484
transform 1 0 31924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_347
timestamp 1666464484
transform 1 0 33028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_359
timestamp 1666464484
transform 1 0 34132 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_366
timestamp 1666464484
transform 1 0 34776 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_378
timestamp 1666464484
transform 1 0 35880 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_390
timestamp 1666464484
transform 1 0 36984 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_402
timestamp 1666464484
transform 1 0 38088 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_409
timestamp 1666464484
transform 1 0 38732 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1666464484
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1666464484
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_445
timestamp 1666464484
transform 1 0 42044 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_452
timestamp 1666464484
transform 1 0 42688 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_464
timestamp 1666464484
transform 1 0 43792 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_476
timestamp 1666464484
transform 1 0 44896 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_488
timestamp 1666464484
transform 1 0 46000 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_495
timestamp 1666464484
transform 1 0 46644 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_507
timestamp 1666464484
transform 1 0 47748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_519
timestamp 1666464484
transform 1 0 48852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_531
timestamp 1666464484
transform 1 0 49956 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_538
timestamp 1666464484
transform 1 0 50600 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_550
timestamp 1666464484
transform 1 0 51704 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_562
timestamp 1666464484
transform 1 0 52808 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_574
timestamp 1666464484
transform 1 0 53912 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_581
timestamp 1666464484
transform 1 0 54556 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_593
timestamp 1666464484
transform 1 0 55660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_605
timestamp 1666464484
transform 1 0 56764 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_617
timestamp 1666464484
transform 1 0 57868 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_624
timestamp 1666464484
transform 1 0 58512 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1666464484
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_39
timestamp 1666464484
transform 1 0 4692 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_44
timestamp 1666464484
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_56
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_68
timestamp 1666464484
transform 1 0 7360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_80
timestamp 1666464484
transform 1 0 8464 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_87
timestamp 1666464484
transform 1 0 9108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_99
timestamp 1666464484
transform 1 0 10212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_123
timestamp 1666464484
transform 1 0 12420 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_130
timestamp 1666464484
transform 1 0 13064 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_142
timestamp 1666464484
transform 1 0 14168 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_154
timestamp 1666464484
transform 1 0 15272 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_166
timestamp 1666464484
transform 1 0 16376 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_173
timestamp 1666464484
transform 1 0 17020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_185
timestamp 1666464484
transform 1 0 18124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_197
timestamp 1666464484
transform 1 0 19228 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_209
timestamp 1666464484
transform 1 0 20332 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_216
timestamp 1666464484
transform 1 0 20976 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_228
timestamp 1666464484
transform 1 0 22080 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_240
timestamp 1666464484
transform 1 0 23184 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_252
timestamp 1666464484
transform 1 0 24288 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_259
timestamp 1666464484
transform 1 0 24932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_271
timestamp 1666464484
transform 1 0 26036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_283
timestamp 1666464484
transform 1 0 27140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_295
timestamp 1666464484
transform 1 0 28244 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_302
timestamp 1666464484
transform 1 0 28888 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_314
timestamp 1666464484
transform 1 0 29992 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_326
timestamp 1666464484
transform 1 0 31096 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_338
timestamp 1666464484
transform 1 0 32200 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_345
timestamp 1666464484
transform 1 0 32844 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_357
timestamp 1666464484
transform 1 0 33948 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_369
timestamp 1666464484
transform 1 0 35052 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_381
timestamp 1666464484
transform 1 0 36156 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_388
timestamp 1666464484
transform 1 0 36800 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_400
timestamp 1666464484
transform 1 0 37904 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_412
timestamp 1666464484
transform 1 0 39008 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_424
timestamp 1666464484
transform 1 0 40112 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_431
timestamp 1666464484
transform 1 0 40756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_443
timestamp 1666464484
transform 1 0 41860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_455
timestamp 1666464484
transform 1 0 42964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_467
timestamp 1666464484
transform 1 0 44068 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_474
timestamp 1666464484
transform 1 0 44712 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_486
timestamp 1666464484
transform 1 0 45816 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_498
timestamp 1666464484
transform 1 0 46920 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_510
timestamp 1666464484
transform 1 0 48024 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1666464484
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1666464484
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1666464484
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1666464484
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_560
timestamp 1666464484
transform 1 0 52624 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_572
timestamp 1666464484
transform 1 0 53728 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_584
timestamp 1666464484
transform 1 0 54832 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_596
timestamp 1666464484
transform 1 0 55936 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_603
timestamp 1666464484
transform 1 0 56580 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_615
timestamp 1666464484
transform 1 0 57684 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_623
timestamp 1666464484
transform 1 0 58420 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_15
timestamp 1666464484
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_22
timestamp 1666464484
transform 1 0 3128 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_34
timestamp 1666464484
transform 1 0 4232 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_46
timestamp 1666464484
transform 1 0 5336 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_58
timestamp 1666464484
transform 1 0 6440 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_89
timestamp 1666464484
transform 1 0 9292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_101
timestamp 1666464484
transform 1 0 10396 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_108
timestamp 1666464484
transform 1 0 11040 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_120
timestamp 1666464484
transform 1 0 12144 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_132
timestamp 1666464484
transform 1 0 13248 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_144
timestamp 1666464484
transform 1 0 14352 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_151
timestamp 1666464484
transform 1 0 14996 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_163
timestamp 1666464484
transform 1 0 16100 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_175
timestamp 1666464484
transform 1 0 17204 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_187
timestamp 1666464484
transform 1 0 18308 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_194
timestamp 1666464484
transform 1 0 18952 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_206
timestamp 1666464484
transform 1 0 20056 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_218
timestamp 1666464484
transform 1 0 21160 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_230
timestamp 1666464484
transform 1 0 22264 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_237
timestamp 1666464484
transform 1 0 22908 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_249
timestamp 1666464484
transform 1 0 24012 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_261
timestamp 1666464484
transform 1 0 25116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_273
timestamp 1666464484
transform 1 0 26220 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_280
timestamp 1666464484
transform 1 0 26864 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_292
timestamp 1666464484
transform 1 0 27968 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_304
timestamp 1666464484
transform 1 0 29072 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_316
timestamp 1666464484
transform 1 0 30176 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_323
timestamp 1666464484
transform 1 0 30820 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_335
timestamp 1666464484
transform 1 0 31924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_347
timestamp 1666464484
transform 1 0 33028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_359
timestamp 1666464484
transform 1 0 34132 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_366
timestamp 1666464484
transform 1 0 34776 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_378
timestamp 1666464484
transform 1 0 35880 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_390
timestamp 1666464484
transform 1 0 36984 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_402
timestamp 1666464484
transform 1 0 38088 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_409
timestamp 1666464484
transform 1 0 38732 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1666464484
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1666464484
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_445
timestamp 1666464484
transform 1 0 42044 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_452
timestamp 1666464484
transform 1 0 42688 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_464
timestamp 1666464484
transform 1 0 43792 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_476
timestamp 1666464484
transform 1 0 44896 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_488
timestamp 1666464484
transform 1 0 46000 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_495
timestamp 1666464484
transform 1 0 46644 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_507
timestamp 1666464484
transform 1 0 47748 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_519
timestamp 1666464484
transform 1 0 48852 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_531
timestamp 1666464484
transform 1 0 49956 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_538
timestamp 1666464484
transform 1 0 50600 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_550
timestamp 1666464484
transform 1 0 51704 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_562
timestamp 1666464484
transform 1 0 52808 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_574
timestamp 1666464484
transform 1 0 53912 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_581
timestamp 1666464484
transform 1 0 54556 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_593
timestamp 1666464484
transform 1 0 55660 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_605
timestamp 1666464484
transform 1 0 56764 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_617
timestamp 1666464484
transform 1 0 57868 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_624
timestamp 1666464484
transform 1 0 58512 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_39
timestamp 1666464484
transform 1 0 4692 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_44
timestamp 1666464484
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_56
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_68
timestamp 1666464484
transform 1 0 7360 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_80
timestamp 1666464484
transform 1 0 8464 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_87
timestamp 1666464484
transform 1 0 9108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_99
timestamp 1666464484
transform 1 0 10212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_123
timestamp 1666464484
transform 1 0 12420 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_130
timestamp 1666464484
transform 1 0 13064 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_142
timestamp 1666464484
transform 1 0 14168 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_154
timestamp 1666464484
transform 1 0 15272 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_166
timestamp 1666464484
transform 1 0 16376 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_173
timestamp 1666464484
transform 1 0 17020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_185
timestamp 1666464484
transform 1 0 18124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_197
timestamp 1666464484
transform 1 0 19228 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_209
timestamp 1666464484
transform 1 0 20332 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_216
timestamp 1666464484
transform 1 0 20976 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_228
timestamp 1666464484
transform 1 0 22080 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_240
timestamp 1666464484
transform 1 0 23184 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_252
timestamp 1666464484
transform 1 0 24288 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_259
timestamp 1666464484
transform 1 0 24932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_271
timestamp 1666464484
transform 1 0 26036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_283
timestamp 1666464484
transform 1 0 27140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_295
timestamp 1666464484
transform 1 0 28244 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_302
timestamp 1666464484
transform 1 0 28888 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_314
timestamp 1666464484
transform 1 0 29992 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_326
timestamp 1666464484
transform 1 0 31096 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_338
timestamp 1666464484
transform 1 0 32200 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_345
timestamp 1666464484
transform 1 0 32844 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_357
timestamp 1666464484
transform 1 0 33948 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_369
timestamp 1666464484
transform 1 0 35052 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_381
timestamp 1666464484
transform 1 0 36156 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_388
timestamp 1666464484
transform 1 0 36800 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_400
timestamp 1666464484
transform 1 0 37904 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_412
timestamp 1666464484
transform 1 0 39008 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_424
timestamp 1666464484
transform 1 0 40112 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_431
timestamp 1666464484
transform 1 0 40756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_443
timestamp 1666464484
transform 1 0 41860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_455
timestamp 1666464484
transform 1 0 42964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_467
timestamp 1666464484
transform 1 0 44068 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_474
timestamp 1666464484
transform 1 0 44712 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_486
timestamp 1666464484
transform 1 0 45816 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_498
timestamp 1666464484
transform 1 0 46920 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_510
timestamp 1666464484
transform 1 0 48024 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1666464484
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1666464484
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1666464484
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1666464484
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_560
timestamp 1666464484
transform 1 0 52624 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_572
timestamp 1666464484
transform 1 0 53728 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_584
timestamp 1666464484
transform 1 0 54832 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_596
timestamp 1666464484
transform 1 0 55936 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_603
timestamp 1666464484
transform 1 0 56580 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_615
timestamp 1666464484
transform 1 0 57684 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_623
timestamp 1666464484
transform 1 0 58420 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_22
timestamp 1666464484
transform 1 0 3128 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_34
timestamp 1666464484
transform 1 0 4232 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_46
timestamp 1666464484
transform 1 0 5336 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_58
timestamp 1666464484
transform 1 0 6440 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_89
timestamp 1666464484
transform 1 0 9292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_101
timestamp 1666464484
transform 1 0 10396 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_108
timestamp 1666464484
transform 1 0 11040 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_120
timestamp 1666464484
transform 1 0 12144 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_132
timestamp 1666464484
transform 1 0 13248 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_144
timestamp 1666464484
transform 1 0 14352 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_151
timestamp 1666464484
transform 1 0 14996 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_163
timestamp 1666464484
transform 1 0 16100 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_175
timestamp 1666464484
transform 1 0 17204 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_187
timestamp 1666464484
transform 1 0 18308 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_194
timestamp 1666464484
transform 1 0 18952 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_206
timestamp 1666464484
transform 1 0 20056 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_218
timestamp 1666464484
transform 1 0 21160 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_230
timestamp 1666464484
transform 1 0 22264 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_237
timestamp 1666464484
transform 1 0 22908 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_249
timestamp 1666464484
transform 1 0 24012 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_261
timestamp 1666464484
transform 1 0 25116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_273
timestamp 1666464484
transform 1 0 26220 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_280
timestamp 1666464484
transform 1 0 26864 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_292
timestamp 1666464484
transform 1 0 27968 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_304
timestamp 1666464484
transform 1 0 29072 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_316
timestamp 1666464484
transform 1 0 30176 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_323
timestamp 1666464484
transform 1 0 30820 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_335
timestamp 1666464484
transform 1 0 31924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_347
timestamp 1666464484
transform 1 0 33028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_359
timestamp 1666464484
transform 1 0 34132 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_366
timestamp 1666464484
transform 1 0 34776 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_378
timestamp 1666464484
transform 1 0 35880 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_390
timestamp 1666464484
transform 1 0 36984 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_402
timestamp 1666464484
transform 1 0 38088 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_409
timestamp 1666464484
transform 1 0 38732 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1666464484
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1666464484
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_445
timestamp 1666464484
transform 1 0 42044 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_452
timestamp 1666464484
transform 1 0 42688 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_464
timestamp 1666464484
transform 1 0 43792 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_476
timestamp 1666464484
transform 1 0 44896 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_488
timestamp 1666464484
transform 1 0 46000 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_495
timestamp 1666464484
transform 1 0 46644 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_507
timestamp 1666464484
transform 1 0 47748 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_519
timestamp 1666464484
transform 1 0 48852 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_531
timestamp 1666464484
transform 1 0 49956 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_538
timestamp 1666464484
transform 1 0 50600 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_550
timestamp 1666464484
transform 1 0 51704 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_562
timestamp 1666464484
transform 1 0 52808 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_574
timestamp 1666464484
transform 1 0 53912 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_581
timestamp 1666464484
transform 1 0 54556 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_593
timestamp 1666464484
transform 1 0 55660 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_605
timestamp 1666464484
transform 1 0 56764 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_617
timestamp 1666464484
transform 1 0 57868 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_624
timestamp 1666464484
transform 1 0 58512 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666464484
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_39
timestamp 1666464484
transform 1 0 4692 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1666464484
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_56
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_68
timestamp 1666464484
transform 1 0 7360 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_80
timestamp 1666464484
transform 1 0 8464 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_87
timestamp 1666464484
transform 1 0 9108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_99
timestamp 1666464484
transform 1 0 10212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_123
timestamp 1666464484
transform 1 0 12420 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_130
timestamp 1666464484
transform 1 0 13064 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_142
timestamp 1666464484
transform 1 0 14168 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_154
timestamp 1666464484
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_166
timestamp 1666464484
transform 1 0 16376 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_173
timestamp 1666464484
transform 1 0 17020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_185
timestamp 1666464484
transform 1 0 18124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_197
timestamp 1666464484
transform 1 0 19228 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_209
timestamp 1666464484
transform 1 0 20332 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_216
timestamp 1666464484
transform 1 0 20976 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_228
timestamp 1666464484
transform 1 0 22080 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_240
timestamp 1666464484
transform 1 0 23184 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_252
timestamp 1666464484
transform 1 0 24288 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_259
timestamp 1666464484
transform 1 0 24932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_271
timestamp 1666464484
transform 1 0 26036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_283
timestamp 1666464484
transform 1 0 27140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_295
timestamp 1666464484
transform 1 0 28244 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_302
timestamp 1666464484
transform 1 0 28888 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_314
timestamp 1666464484
transform 1 0 29992 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_326
timestamp 1666464484
transform 1 0 31096 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_338
timestamp 1666464484
transform 1 0 32200 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_345
timestamp 1666464484
transform 1 0 32844 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_357
timestamp 1666464484
transform 1 0 33948 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_369
timestamp 1666464484
transform 1 0 35052 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_381
timestamp 1666464484
transform 1 0 36156 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_388
timestamp 1666464484
transform 1 0 36800 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_400
timestamp 1666464484
transform 1 0 37904 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_412
timestamp 1666464484
transform 1 0 39008 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_424
timestamp 1666464484
transform 1 0 40112 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_431
timestamp 1666464484
transform 1 0 40756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_443
timestamp 1666464484
transform 1 0 41860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_455
timestamp 1666464484
transform 1 0 42964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_467
timestamp 1666464484
transform 1 0 44068 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_474
timestamp 1666464484
transform 1 0 44712 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_486
timestamp 1666464484
transform 1 0 45816 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_498
timestamp 1666464484
transform 1 0 46920 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_510
timestamp 1666464484
transform 1 0 48024 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1666464484
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1666464484
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1666464484
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1666464484
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_560
timestamp 1666464484
transform 1 0 52624 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_572
timestamp 1666464484
transform 1 0 53728 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_584
timestamp 1666464484
transform 1 0 54832 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_596
timestamp 1666464484
transform 1 0 55936 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_603
timestamp 1666464484
transform 1 0 56580 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_615
timestamp 1666464484
transform 1 0 57684 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_623
timestamp 1666464484
transform 1 0 58420 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_22
timestamp 1666464484
transform 1 0 3128 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_34
timestamp 1666464484
transform 1 0 4232 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_46
timestamp 1666464484
transform 1 0 5336 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_58
timestamp 1666464484
transform 1 0 6440 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_89
timestamp 1666464484
transform 1 0 9292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_101
timestamp 1666464484
transform 1 0 10396 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_108
timestamp 1666464484
transform 1 0 11040 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_120
timestamp 1666464484
transform 1 0 12144 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_132
timestamp 1666464484
transform 1 0 13248 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_144
timestamp 1666464484
transform 1 0 14352 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_151
timestamp 1666464484
transform 1 0 14996 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_163
timestamp 1666464484
transform 1 0 16100 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_175
timestamp 1666464484
transform 1 0 17204 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_187
timestamp 1666464484
transform 1 0 18308 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_194
timestamp 1666464484
transform 1 0 18952 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_206
timestamp 1666464484
transform 1 0 20056 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_218
timestamp 1666464484
transform 1 0 21160 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_230
timestamp 1666464484
transform 1 0 22264 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_237
timestamp 1666464484
transform 1 0 22908 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_249
timestamp 1666464484
transform 1 0 24012 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_261
timestamp 1666464484
transform 1 0 25116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_273
timestamp 1666464484
transform 1 0 26220 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_280
timestamp 1666464484
transform 1 0 26864 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_292
timestamp 1666464484
transform 1 0 27968 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_304
timestamp 1666464484
transform 1 0 29072 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_316
timestamp 1666464484
transform 1 0 30176 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_323
timestamp 1666464484
transform 1 0 30820 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_335
timestamp 1666464484
transform 1 0 31924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_347
timestamp 1666464484
transform 1 0 33028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_359
timestamp 1666464484
transform 1 0 34132 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_366
timestamp 1666464484
transform 1 0 34776 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_378
timestamp 1666464484
transform 1 0 35880 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_390
timestamp 1666464484
transform 1 0 36984 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_402
timestamp 1666464484
transform 1 0 38088 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_409
timestamp 1666464484
transform 1 0 38732 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1666464484
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1666464484
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_445
timestamp 1666464484
transform 1 0 42044 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_452
timestamp 1666464484
transform 1 0 42688 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_464
timestamp 1666464484
transform 1 0 43792 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_476
timestamp 1666464484
transform 1 0 44896 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_488
timestamp 1666464484
transform 1 0 46000 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_495
timestamp 1666464484
transform 1 0 46644 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_507
timestamp 1666464484
transform 1 0 47748 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_519
timestamp 1666464484
transform 1 0 48852 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_531
timestamp 1666464484
transform 1 0 49956 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_538
timestamp 1666464484
transform 1 0 50600 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_550
timestamp 1666464484
transform 1 0 51704 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_562
timestamp 1666464484
transform 1 0 52808 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_574
timestamp 1666464484
transform 1 0 53912 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_581
timestamp 1666464484
transform 1 0 54556 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_593
timestamp 1666464484
transform 1 0 55660 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_605
timestamp 1666464484
transform 1 0 56764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_617
timestamp 1666464484
transform 1 0 57868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_624
timestamp 1666464484
transform 1 0 58512 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_44
timestamp 1666464484
transform 1 0 5152 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_56
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_68
timestamp 1666464484
transform 1 0 7360 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_80
timestamp 1666464484
transform 1 0 8464 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_87
timestamp 1666464484
transform 1 0 9108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_99
timestamp 1666464484
transform 1 0 10212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_123
timestamp 1666464484
transform 1 0 12420 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_130
timestamp 1666464484
transform 1 0 13064 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_142
timestamp 1666464484
transform 1 0 14168 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_154
timestamp 1666464484
transform 1 0 15272 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_166
timestamp 1666464484
transform 1 0 16376 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_173
timestamp 1666464484
transform 1 0 17020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_185
timestamp 1666464484
transform 1 0 18124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_197
timestamp 1666464484
transform 1 0 19228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_209
timestamp 1666464484
transform 1 0 20332 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_216
timestamp 1666464484
transform 1 0 20976 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_228
timestamp 1666464484
transform 1 0 22080 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_240
timestamp 1666464484
transform 1 0 23184 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_252
timestamp 1666464484
transform 1 0 24288 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_259
timestamp 1666464484
transform 1 0 24932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_271
timestamp 1666464484
transform 1 0 26036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_283
timestamp 1666464484
transform 1 0 27140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_295
timestamp 1666464484
transform 1 0 28244 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_302
timestamp 1666464484
transform 1 0 28888 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_314
timestamp 1666464484
transform 1 0 29992 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_326
timestamp 1666464484
transform 1 0 31096 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_338
timestamp 1666464484
transform 1 0 32200 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_345
timestamp 1666464484
transform 1 0 32844 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_357
timestamp 1666464484
transform 1 0 33948 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_369
timestamp 1666464484
transform 1 0 35052 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_381
timestamp 1666464484
transform 1 0 36156 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_388
timestamp 1666464484
transform 1 0 36800 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_400
timestamp 1666464484
transform 1 0 37904 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_412
timestamp 1666464484
transform 1 0 39008 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_424
timestamp 1666464484
transform 1 0 40112 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_431
timestamp 1666464484
transform 1 0 40756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_443
timestamp 1666464484
transform 1 0 41860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_455
timestamp 1666464484
transform 1 0 42964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_467
timestamp 1666464484
transform 1 0 44068 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_474
timestamp 1666464484
transform 1 0 44712 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_486
timestamp 1666464484
transform 1 0 45816 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_498
timestamp 1666464484
transform 1 0 46920 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_510
timestamp 1666464484
transform 1 0 48024 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1666464484
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1666464484
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1666464484
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1666464484
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_560
timestamp 1666464484
transform 1 0 52624 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_572
timestamp 1666464484
transform 1 0 53728 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_584
timestamp 1666464484
transform 1 0 54832 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_596
timestamp 1666464484
transform 1 0 55936 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_603
timestamp 1666464484
transform 1 0 56580 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_615
timestamp 1666464484
transform 1 0 57684 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_623
timestamp 1666464484
transform 1 0 58420 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_15
timestamp 1666464484
transform 1 0 2484 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_22
timestamp 1666464484
transform 1 0 3128 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_34
timestamp 1666464484
transform 1 0 4232 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_46
timestamp 1666464484
transform 1 0 5336 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_58
timestamp 1666464484
transform 1 0 6440 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_89
timestamp 1666464484
transform 1 0 9292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_101
timestamp 1666464484
transform 1 0 10396 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_108
timestamp 1666464484
transform 1 0 11040 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_120
timestamp 1666464484
transform 1 0 12144 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_132
timestamp 1666464484
transform 1 0 13248 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_144
timestamp 1666464484
transform 1 0 14352 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_151
timestamp 1666464484
transform 1 0 14996 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_163
timestamp 1666464484
transform 1 0 16100 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_175
timestamp 1666464484
transform 1 0 17204 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_187
timestamp 1666464484
transform 1 0 18308 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_194
timestamp 1666464484
transform 1 0 18952 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_206
timestamp 1666464484
transform 1 0 20056 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_218
timestamp 1666464484
transform 1 0 21160 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_230
timestamp 1666464484
transform 1 0 22264 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_237
timestamp 1666464484
transform 1 0 22908 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_249
timestamp 1666464484
transform 1 0 24012 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_261
timestamp 1666464484
transform 1 0 25116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_273
timestamp 1666464484
transform 1 0 26220 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_280
timestamp 1666464484
transform 1 0 26864 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_292
timestamp 1666464484
transform 1 0 27968 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_304
timestamp 1666464484
transform 1 0 29072 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_316
timestamp 1666464484
transform 1 0 30176 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_323
timestamp 1666464484
transform 1 0 30820 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_335
timestamp 1666464484
transform 1 0 31924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_347
timestamp 1666464484
transform 1 0 33028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_359
timestamp 1666464484
transform 1 0 34132 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_366
timestamp 1666464484
transform 1 0 34776 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_378
timestamp 1666464484
transform 1 0 35880 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_390
timestamp 1666464484
transform 1 0 36984 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_402
timestamp 1666464484
transform 1 0 38088 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_409
timestamp 1666464484
transform 1 0 38732 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1666464484
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1666464484
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_445
timestamp 1666464484
transform 1 0 42044 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_452
timestamp 1666464484
transform 1 0 42688 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_464
timestamp 1666464484
transform 1 0 43792 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_476
timestamp 1666464484
transform 1 0 44896 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_488
timestamp 1666464484
transform 1 0 46000 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_495
timestamp 1666464484
transform 1 0 46644 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_507
timestamp 1666464484
transform 1 0 47748 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_519
timestamp 1666464484
transform 1 0 48852 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_531
timestamp 1666464484
transform 1 0 49956 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_538
timestamp 1666464484
transform 1 0 50600 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_550
timestamp 1666464484
transform 1 0 51704 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_562
timestamp 1666464484
transform 1 0 52808 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_574
timestamp 1666464484
transform 1 0 53912 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_581
timestamp 1666464484
transform 1 0 54556 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_593
timestamp 1666464484
transform 1 0 55660 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_605
timestamp 1666464484
transform 1 0 56764 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_617
timestamp 1666464484
transform 1 0 57868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_624
timestamp 1666464484
transform 1 0 58512 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_44
timestamp 1666464484
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_56
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_68
timestamp 1666464484
transform 1 0 7360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_80
timestamp 1666464484
transform 1 0 8464 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_87
timestamp 1666464484
transform 1 0 9108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_99
timestamp 1666464484
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_123
timestamp 1666464484
transform 1 0 12420 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_130
timestamp 1666464484
transform 1 0 13064 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_142
timestamp 1666464484
transform 1 0 14168 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_154
timestamp 1666464484
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_166
timestamp 1666464484
transform 1 0 16376 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_173
timestamp 1666464484
transform 1 0 17020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_185
timestamp 1666464484
transform 1 0 18124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_197
timestamp 1666464484
transform 1 0 19228 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_209
timestamp 1666464484
transform 1 0 20332 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_216
timestamp 1666464484
transform 1 0 20976 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_228
timestamp 1666464484
transform 1 0 22080 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_240
timestamp 1666464484
transform 1 0 23184 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_252
timestamp 1666464484
transform 1 0 24288 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_259
timestamp 1666464484
transform 1 0 24932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_271
timestamp 1666464484
transform 1 0 26036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_283
timestamp 1666464484
transform 1 0 27140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_295
timestamp 1666464484
transform 1 0 28244 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_302
timestamp 1666464484
transform 1 0 28888 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_314
timestamp 1666464484
transform 1 0 29992 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_326
timestamp 1666464484
transform 1 0 31096 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_338
timestamp 1666464484
transform 1 0 32200 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_345
timestamp 1666464484
transform 1 0 32844 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_357
timestamp 1666464484
transform 1 0 33948 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_369
timestamp 1666464484
transform 1 0 35052 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_381
timestamp 1666464484
transform 1 0 36156 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_388
timestamp 1666464484
transform 1 0 36800 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_400
timestamp 1666464484
transform 1 0 37904 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_412
timestamp 1666464484
transform 1 0 39008 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_424
timestamp 1666464484
transform 1 0 40112 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_431
timestamp 1666464484
transform 1 0 40756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_443
timestamp 1666464484
transform 1 0 41860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_455
timestamp 1666464484
transform 1 0 42964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_467
timestamp 1666464484
transform 1 0 44068 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_474
timestamp 1666464484
transform 1 0 44712 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_486
timestamp 1666464484
transform 1 0 45816 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_498
timestamp 1666464484
transform 1 0 46920 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_510
timestamp 1666464484
transform 1 0 48024 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1666464484
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1666464484
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1666464484
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1666464484
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_560
timestamp 1666464484
transform 1 0 52624 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_572
timestamp 1666464484
transform 1 0 53728 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_584
timestamp 1666464484
transform 1 0 54832 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_596
timestamp 1666464484
transform 1 0 55936 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_603
timestamp 1666464484
transform 1 0 56580 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_615
timestamp 1666464484
transform 1 0 57684 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_623
timestamp 1666464484
transform 1 0 58420 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_15
timestamp 1666464484
transform 1 0 2484 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_22
timestamp 1666464484
transform 1 0 3128 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_34
timestamp 1666464484
transform 1 0 4232 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_46
timestamp 1666464484
transform 1 0 5336 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_58
timestamp 1666464484
transform 1 0 6440 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_89
timestamp 1666464484
transform 1 0 9292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_101
timestamp 1666464484
transform 1 0 10396 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_108
timestamp 1666464484
transform 1 0 11040 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_120
timestamp 1666464484
transform 1 0 12144 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_132
timestamp 1666464484
transform 1 0 13248 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_144
timestamp 1666464484
transform 1 0 14352 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_151
timestamp 1666464484
transform 1 0 14996 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_163
timestamp 1666464484
transform 1 0 16100 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_175
timestamp 1666464484
transform 1 0 17204 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_187
timestamp 1666464484
transform 1 0 18308 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_194
timestamp 1666464484
transform 1 0 18952 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_206
timestamp 1666464484
transform 1 0 20056 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_218
timestamp 1666464484
transform 1 0 21160 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_230
timestamp 1666464484
transform 1 0 22264 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_237
timestamp 1666464484
transform 1 0 22908 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_249
timestamp 1666464484
transform 1 0 24012 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_261
timestamp 1666464484
transform 1 0 25116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_273
timestamp 1666464484
transform 1 0 26220 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_280
timestamp 1666464484
transform 1 0 26864 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_292
timestamp 1666464484
transform 1 0 27968 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_304
timestamp 1666464484
transform 1 0 29072 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_316
timestamp 1666464484
transform 1 0 30176 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_323
timestamp 1666464484
transform 1 0 30820 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_335
timestamp 1666464484
transform 1 0 31924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_347
timestamp 1666464484
transform 1 0 33028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_359
timestamp 1666464484
transform 1 0 34132 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_366
timestamp 1666464484
transform 1 0 34776 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_378
timestamp 1666464484
transform 1 0 35880 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_390
timestamp 1666464484
transform 1 0 36984 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_402
timestamp 1666464484
transform 1 0 38088 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_409
timestamp 1666464484
transform 1 0 38732 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1666464484
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1666464484
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_445
timestamp 1666464484
transform 1 0 42044 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_452
timestamp 1666464484
transform 1 0 42688 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_464
timestamp 1666464484
transform 1 0 43792 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_476
timestamp 1666464484
transform 1 0 44896 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_488
timestamp 1666464484
transform 1 0 46000 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_495
timestamp 1666464484
transform 1 0 46644 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_507
timestamp 1666464484
transform 1 0 47748 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_519
timestamp 1666464484
transform 1 0 48852 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_531
timestamp 1666464484
transform 1 0 49956 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_538
timestamp 1666464484
transform 1 0 50600 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_550
timestamp 1666464484
transform 1 0 51704 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_562
timestamp 1666464484
transform 1 0 52808 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_574
timestamp 1666464484
transform 1 0 53912 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_581
timestamp 1666464484
transform 1 0 54556 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_593
timestamp 1666464484
transform 1 0 55660 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_605
timestamp 1666464484
transform 1 0 56764 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_617
timestamp 1666464484
transform 1 0 57868 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_624
timestamp 1666464484
transform 1 0 58512 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_39
timestamp 1666464484
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_44
timestamp 1666464484
transform 1 0 5152 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_56
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_68
timestamp 1666464484
transform 1 0 7360 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_80
timestamp 1666464484
transform 1 0 8464 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_87
timestamp 1666464484
transform 1 0 9108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_99
timestamp 1666464484
transform 1 0 10212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_123
timestamp 1666464484
transform 1 0 12420 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_130
timestamp 1666464484
transform 1 0 13064 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_142
timestamp 1666464484
transform 1 0 14168 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_154
timestamp 1666464484
transform 1 0 15272 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_166
timestamp 1666464484
transform 1 0 16376 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_173
timestamp 1666464484
transform 1 0 17020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_185
timestamp 1666464484
transform 1 0 18124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_197
timestamp 1666464484
transform 1 0 19228 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_209
timestamp 1666464484
transform 1 0 20332 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_216
timestamp 1666464484
transform 1 0 20976 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_228
timestamp 1666464484
transform 1 0 22080 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_240
timestamp 1666464484
transform 1 0 23184 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_252
timestamp 1666464484
transform 1 0 24288 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_259
timestamp 1666464484
transform 1 0 24932 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_271
timestamp 1666464484
transform 1 0 26036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_283
timestamp 1666464484
transform 1 0 27140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_295
timestamp 1666464484
transform 1 0 28244 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_302
timestamp 1666464484
transform 1 0 28888 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_314
timestamp 1666464484
transform 1 0 29992 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_326
timestamp 1666464484
transform 1 0 31096 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_338
timestamp 1666464484
transform 1 0 32200 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_345
timestamp 1666464484
transform 1 0 32844 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_357
timestamp 1666464484
transform 1 0 33948 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_369
timestamp 1666464484
transform 1 0 35052 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_381
timestamp 1666464484
transform 1 0 36156 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_388
timestamp 1666464484
transform 1 0 36800 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_400
timestamp 1666464484
transform 1 0 37904 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_412
timestamp 1666464484
transform 1 0 39008 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_424
timestamp 1666464484
transform 1 0 40112 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_431
timestamp 1666464484
transform 1 0 40756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_443
timestamp 1666464484
transform 1 0 41860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_455
timestamp 1666464484
transform 1 0 42964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_467
timestamp 1666464484
transform 1 0 44068 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_474
timestamp 1666464484
transform 1 0 44712 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_486
timestamp 1666464484
transform 1 0 45816 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_498
timestamp 1666464484
transform 1 0 46920 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_510
timestamp 1666464484
transform 1 0 48024 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1666464484
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1666464484
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1666464484
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1666464484
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_560
timestamp 1666464484
transform 1 0 52624 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_572
timestamp 1666464484
transform 1 0 53728 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_584
timestamp 1666464484
transform 1 0 54832 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_596
timestamp 1666464484
transform 1 0 55936 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_603
timestamp 1666464484
transform 1 0 56580 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_615
timestamp 1666464484
transform 1 0 57684 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_623
timestamp 1666464484
transform 1 0 58420 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_22
timestamp 1666464484
transform 1 0 3128 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_34
timestamp 1666464484
transform 1 0 4232 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_46
timestamp 1666464484
transform 1 0 5336 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_58
timestamp 1666464484
transform 1 0 6440 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_89
timestamp 1666464484
transform 1 0 9292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_101
timestamp 1666464484
transform 1 0 10396 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_108
timestamp 1666464484
transform 1 0 11040 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_120
timestamp 1666464484
transform 1 0 12144 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_132
timestamp 1666464484
transform 1 0 13248 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_144
timestamp 1666464484
transform 1 0 14352 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_151
timestamp 1666464484
transform 1 0 14996 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_163
timestamp 1666464484
transform 1 0 16100 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_175
timestamp 1666464484
transform 1 0 17204 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_187
timestamp 1666464484
transform 1 0 18308 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_194
timestamp 1666464484
transform 1 0 18952 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_206
timestamp 1666464484
transform 1 0 20056 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_218
timestamp 1666464484
transform 1 0 21160 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_230
timestamp 1666464484
transform 1 0 22264 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_237
timestamp 1666464484
transform 1 0 22908 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_249
timestamp 1666464484
transform 1 0 24012 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_261
timestamp 1666464484
transform 1 0 25116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_273
timestamp 1666464484
transform 1 0 26220 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_280
timestamp 1666464484
transform 1 0 26864 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_292
timestamp 1666464484
transform 1 0 27968 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_304
timestamp 1666464484
transform 1 0 29072 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_316
timestamp 1666464484
transform 1 0 30176 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_323
timestamp 1666464484
transform 1 0 30820 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_335
timestamp 1666464484
transform 1 0 31924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_347
timestamp 1666464484
transform 1 0 33028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_359
timestamp 1666464484
transform 1 0 34132 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_366
timestamp 1666464484
transform 1 0 34776 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_378
timestamp 1666464484
transform 1 0 35880 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_390
timestamp 1666464484
transform 1 0 36984 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_402
timestamp 1666464484
transform 1 0 38088 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_409
timestamp 1666464484
transform 1 0 38732 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1666464484
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1666464484
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_445
timestamp 1666464484
transform 1 0 42044 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_452
timestamp 1666464484
transform 1 0 42688 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_464
timestamp 1666464484
transform 1 0 43792 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_476
timestamp 1666464484
transform 1 0 44896 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_488
timestamp 1666464484
transform 1 0 46000 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_495
timestamp 1666464484
transform 1 0 46644 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_507
timestamp 1666464484
transform 1 0 47748 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_519
timestamp 1666464484
transform 1 0 48852 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_531
timestamp 1666464484
transform 1 0 49956 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_538
timestamp 1666464484
transform 1 0 50600 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_550
timestamp 1666464484
transform 1 0 51704 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_562
timestamp 1666464484
transform 1 0 52808 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_574
timestamp 1666464484
transform 1 0 53912 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_581
timestamp 1666464484
transform 1 0 54556 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_593
timestamp 1666464484
transform 1 0 55660 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_605
timestamp 1666464484
transform 1 0 56764 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_617
timestamp 1666464484
transform 1 0 57868 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_624
timestamp 1666464484
transform 1 0 58512 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_39
timestamp 1666464484
transform 1 0 4692 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_44
timestamp 1666464484
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_56
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_68
timestamp 1666464484
transform 1 0 7360 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_80
timestamp 1666464484
transform 1 0 8464 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_87
timestamp 1666464484
transform 1 0 9108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_99
timestamp 1666464484
transform 1 0 10212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_123
timestamp 1666464484
transform 1 0 12420 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_130
timestamp 1666464484
transform 1 0 13064 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_142
timestamp 1666464484
transform 1 0 14168 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_154
timestamp 1666464484
transform 1 0 15272 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_166
timestamp 1666464484
transform 1 0 16376 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_173
timestamp 1666464484
transform 1 0 17020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_185
timestamp 1666464484
transform 1 0 18124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_197
timestamp 1666464484
transform 1 0 19228 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_209
timestamp 1666464484
transform 1 0 20332 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_216
timestamp 1666464484
transform 1 0 20976 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_228
timestamp 1666464484
transform 1 0 22080 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_240
timestamp 1666464484
transform 1 0 23184 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_252
timestamp 1666464484
transform 1 0 24288 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_259
timestamp 1666464484
transform 1 0 24932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_271
timestamp 1666464484
transform 1 0 26036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_283
timestamp 1666464484
transform 1 0 27140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_295
timestamp 1666464484
transform 1 0 28244 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_302
timestamp 1666464484
transform 1 0 28888 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_314
timestamp 1666464484
transform 1 0 29992 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_326
timestamp 1666464484
transform 1 0 31096 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_338
timestamp 1666464484
transform 1 0 32200 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_345
timestamp 1666464484
transform 1 0 32844 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_357
timestamp 1666464484
transform 1 0 33948 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_369
timestamp 1666464484
transform 1 0 35052 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_381
timestamp 1666464484
transform 1 0 36156 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_388
timestamp 1666464484
transform 1 0 36800 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_400
timestamp 1666464484
transform 1 0 37904 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_412
timestamp 1666464484
transform 1 0 39008 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_424
timestamp 1666464484
transform 1 0 40112 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_431
timestamp 1666464484
transform 1 0 40756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_443
timestamp 1666464484
transform 1 0 41860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_455
timestamp 1666464484
transform 1 0 42964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_467
timestamp 1666464484
transform 1 0 44068 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_474
timestamp 1666464484
transform 1 0 44712 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_486
timestamp 1666464484
transform 1 0 45816 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_498
timestamp 1666464484
transform 1 0 46920 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_510
timestamp 1666464484
transform 1 0 48024 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1666464484
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1666464484
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1666464484
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1666464484
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_560
timestamp 1666464484
transform 1 0 52624 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_572
timestamp 1666464484
transform 1 0 53728 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_584
timestamp 1666464484
transform 1 0 54832 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_596
timestamp 1666464484
transform 1 0 55936 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_603
timestamp 1666464484
transform 1 0 56580 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_615
timestamp 1666464484
transform 1 0 57684 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_623
timestamp 1666464484
transform 1 0 58420 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_22
timestamp 1666464484
transform 1 0 3128 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_34
timestamp 1666464484
transform 1 0 4232 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_46
timestamp 1666464484
transform 1 0 5336 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_58
timestamp 1666464484
transform 1 0 6440 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_89
timestamp 1666464484
transform 1 0 9292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_101
timestamp 1666464484
transform 1 0 10396 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_108
timestamp 1666464484
transform 1 0 11040 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_120
timestamp 1666464484
transform 1 0 12144 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_132
timestamp 1666464484
transform 1 0 13248 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_144
timestamp 1666464484
transform 1 0 14352 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_151
timestamp 1666464484
transform 1 0 14996 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_163
timestamp 1666464484
transform 1 0 16100 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_175
timestamp 1666464484
transform 1 0 17204 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_187
timestamp 1666464484
transform 1 0 18308 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_194
timestamp 1666464484
transform 1 0 18952 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_206
timestamp 1666464484
transform 1 0 20056 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_218
timestamp 1666464484
transform 1 0 21160 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_230
timestamp 1666464484
transform 1 0 22264 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_237
timestamp 1666464484
transform 1 0 22908 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_249
timestamp 1666464484
transform 1 0 24012 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_261
timestamp 1666464484
transform 1 0 25116 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_273
timestamp 1666464484
transform 1 0 26220 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_280
timestamp 1666464484
transform 1 0 26864 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_292
timestamp 1666464484
transform 1 0 27968 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_304
timestamp 1666464484
transform 1 0 29072 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_316
timestamp 1666464484
transform 1 0 30176 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_323
timestamp 1666464484
transform 1 0 30820 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_335
timestamp 1666464484
transform 1 0 31924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_347
timestamp 1666464484
transform 1 0 33028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_359
timestamp 1666464484
transform 1 0 34132 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_366
timestamp 1666464484
transform 1 0 34776 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_378
timestamp 1666464484
transform 1 0 35880 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_390
timestamp 1666464484
transform 1 0 36984 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_402
timestamp 1666464484
transform 1 0 38088 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_409
timestamp 1666464484
transform 1 0 38732 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1666464484
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1666464484
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_445
timestamp 1666464484
transform 1 0 42044 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_452
timestamp 1666464484
transform 1 0 42688 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_464
timestamp 1666464484
transform 1 0 43792 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_476
timestamp 1666464484
transform 1 0 44896 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_488
timestamp 1666464484
transform 1 0 46000 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_495
timestamp 1666464484
transform 1 0 46644 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_507
timestamp 1666464484
transform 1 0 47748 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_519
timestamp 1666464484
transform 1 0 48852 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_531
timestamp 1666464484
transform 1 0 49956 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_538
timestamp 1666464484
transform 1 0 50600 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_550
timestamp 1666464484
transform 1 0 51704 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_562
timestamp 1666464484
transform 1 0 52808 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_574
timestamp 1666464484
transform 1 0 53912 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_581
timestamp 1666464484
transform 1 0 54556 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_593
timestamp 1666464484
transform 1 0 55660 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_605
timestamp 1666464484
transform 1 0 56764 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_617
timestamp 1666464484
transform 1 0 57868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_624
timestamp 1666464484
transform 1 0 58512 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_44
timestamp 1666464484
transform 1 0 5152 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_56
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_68
timestamp 1666464484
transform 1 0 7360 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_80
timestamp 1666464484
transform 1 0 8464 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_87
timestamp 1666464484
transform 1 0 9108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_99
timestamp 1666464484
transform 1 0 10212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_123
timestamp 1666464484
transform 1 0 12420 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_130
timestamp 1666464484
transform 1 0 13064 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_142
timestamp 1666464484
transform 1 0 14168 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_154
timestamp 1666464484
transform 1 0 15272 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_166
timestamp 1666464484
transform 1 0 16376 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_173
timestamp 1666464484
transform 1 0 17020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_185
timestamp 1666464484
transform 1 0 18124 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_197
timestamp 1666464484
transform 1 0 19228 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_209
timestamp 1666464484
transform 1 0 20332 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_216
timestamp 1666464484
transform 1 0 20976 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_228
timestamp 1666464484
transform 1 0 22080 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_240
timestamp 1666464484
transform 1 0 23184 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_252
timestamp 1666464484
transform 1 0 24288 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_259
timestamp 1666464484
transform 1 0 24932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_271
timestamp 1666464484
transform 1 0 26036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_283
timestamp 1666464484
transform 1 0 27140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_295
timestamp 1666464484
transform 1 0 28244 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_302
timestamp 1666464484
transform 1 0 28888 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_314
timestamp 1666464484
transform 1 0 29992 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_326
timestamp 1666464484
transform 1 0 31096 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_338
timestamp 1666464484
transform 1 0 32200 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_345
timestamp 1666464484
transform 1 0 32844 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_357
timestamp 1666464484
transform 1 0 33948 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_369
timestamp 1666464484
transform 1 0 35052 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_381
timestamp 1666464484
transform 1 0 36156 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_388
timestamp 1666464484
transform 1 0 36800 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_400
timestamp 1666464484
transform 1 0 37904 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_412
timestamp 1666464484
transform 1 0 39008 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_424
timestamp 1666464484
transform 1 0 40112 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_431
timestamp 1666464484
transform 1 0 40756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_443
timestamp 1666464484
transform 1 0 41860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_455
timestamp 1666464484
transform 1 0 42964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_467
timestamp 1666464484
transform 1 0 44068 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_474
timestamp 1666464484
transform 1 0 44712 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_486
timestamp 1666464484
transform 1 0 45816 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_498
timestamp 1666464484
transform 1 0 46920 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_510
timestamp 1666464484
transform 1 0 48024 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1666464484
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1666464484
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1666464484
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1666464484
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_560
timestamp 1666464484
transform 1 0 52624 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_572
timestamp 1666464484
transform 1 0 53728 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_584
timestamp 1666464484
transform 1 0 54832 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_596
timestamp 1666464484
transform 1 0 55936 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_603
timestamp 1666464484
transform 1 0 56580 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_615
timestamp 1666464484
transform 1 0 57684 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_623
timestamp 1666464484
transform 1 0 58420 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_15
timestamp 1666464484
transform 1 0 2484 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_22
timestamp 1666464484
transform 1 0 3128 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_34
timestamp 1666464484
transform 1 0 4232 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_46
timestamp 1666464484
transform 1 0 5336 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_58
timestamp 1666464484
transform 1 0 6440 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_89
timestamp 1666464484
transform 1 0 9292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_101
timestamp 1666464484
transform 1 0 10396 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_108
timestamp 1666464484
transform 1 0 11040 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_120
timestamp 1666464484
transform 1 0 12144 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_132
timestamp 1666464484
transform 1 0 13248 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_144
timestamp 1666464484
transform 1 0 14352 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_151
timestamp 1666464484
transform 1 0 14996 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_163
timestamp 1666464484
transform 1 0 16100 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_175
timestamp 1666464484
transform 1 0 17204 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_187
timestamp 1666464484
transform 1 0 18308 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_194
timestamp 1666464484
transform 1 0 18952 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_206
timestamp 1666464484
transform 1 0 20056 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_218
timestamp 1666464484
transform 1 0 21160 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_230
timestamp 1666464484
transform 1 0 22264 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_237
timestamp 1666464484
transform 1 0 22908 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_249
timestamp 1666464484
transform 1 0 24012 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_261
timestamp 1666464484
transform 1 0 25116 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_273
timestamp 1666464484
transform 1 0 26220 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_280
timestamp 1666464484
transform 1 0 26864 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_292
timestamp 1666464484
transform 1 0 27968 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_304
timestamp 1666464484
transform 1 0 29072 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_316
timestamp 1666464484
transform 1 0 30176 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_323
timestamp 1666464484
transform 1 0 30820 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_335
timestamp 1666464484
transform 1 0 31924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_347
timestamp 1666464484
transform 1 0 33028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_359
timestamp 1666464484
transform 1 0 34132 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_366
timestamp 1666464484
transform 1 0 34776 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_378
timestamp 1666464484
transform 1 0 35880 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_390
timestamp 1666464484
transform 1 0 36984 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_402
timestamp 1666464484
transform 1 0 38088 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_409
timestamp 1666464484
transform 1 0 38732 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1666464484
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1666464484
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_445
timestamp 1666464484
transform 1 0 42044 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_452
timestamp 1666464484
transform 1 0 42688 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_464
timestamp 1666464484
transform 1 0 43792 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_476
timestamp 1666464484
transform 1 0 44896 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_488
timestamp 1666464484
transform 1 0 46000 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_495
timestamp 1666464484
transform 1 0 46644 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_507
timestamp 1666464484
transform 1 0 47748 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_519
timestamp 1666464484
transform 1 0 48852 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_531
timestamp 1666464484
transform 1 0 49956 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_538
timestamp 1666464484
transform 1 0 50600 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_550
timestamp 1666464484
transform 1 0 51704 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_562
timestamp 1666464484
transform 1 0 52808 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_574
timestamp 1666464484
transform 1 0 53912 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_581
timestamp 1666464484
transform 1 0 54556 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_593
timestamp 1666464484
transform 1 0 55660 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_605
timestamp 1666464484
transform 1 0 56764 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_617
timestamp 1666464484
transform 1 0 57868 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_624
timestamp 1666464484
transform 1 0 58512 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666464484
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1666464484
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_39
timestamp 1666464484
transform 1 0 4692 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1666464484
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_56
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_68
timestamp 1666464484
transform 1 0 7360 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_80
timestamp 1666464484
transform 1 0 8464 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_87
timestamp 1666464484
transform 1 0 9108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_99
timestamp 1666464484
transform 1 0 10212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_123
timestamp 1666464484
transform 1 0 12420 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_130
timestamp 1666464484
transform 1 0 13064 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_142
timestamp 1666464484
transform 1 0 14168 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_154
timestamp 1666464484
transform 1 0 15272 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_166
timestamp 1666464484
transform 1 0 16376 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_173
timestamp 1666464484
transform 1 0 17020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_185
timestamp 1666464484
transform 1 0 18124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_197
timestamp 1666464484
transform 1 0 19228 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_209
timestamp 1666464484
transform 1 0 20332 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_216
timestamp 1666464484
transform 1 0 20976 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_228
timestamp 1666464484
transform 1 0 22080 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_240
timestamp 1666464484
transform 1 0 23184 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_252
timestamp 1666464484
transform 1 0 24288 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_259
timestamp 1666464484
transform 1 0 24932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_271
timestamp 1666464484
transform 1 0 26036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_283
timestamp 1666464484
transform 1 0 27140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_295
timestamp 1666464484
transform 1 0 28244 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_302
timestamp 1666464484
transform 1 0 28888 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_314
timestamp 1666464484
transform 1 0 29992 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_326
timestamp 1666464484
transform 1 0 31096 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_338
timestamp 1666464484
transform 1 0 32200 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_345
timestamp 1666464484
transform 1 0 32844 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_357
timestamp 1666464484
transform 1 0 33948 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_369
timestamp 1666464484
transform 1 0 35052 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_381
timestamp 1666464484
transform 1 0 36156 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_388
timestamp 1666464484
transform 1 0 36800 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_400
timestamp 1666464484
transform 1 0 37904 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_412
timestamp 1666464484
transform 1 0 39008 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_424
timestamp 1666464484
transform 1 0 40112 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_431
timestamp 1666464484
transform 1 0 40756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_443
timestamp 1666464484
transform 1 0 41860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_455
timestamp 1666464484
transform 1 0 42964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_467
timestamp 1666464484
transform 1 0 44068 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_474
timestamp 1666464484
transform 1 0 44712 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_486
timestamp 1666464484
transform 1 0 45816 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_498
timestamp 1666464484
transform 1 0 46920 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_510
timestamp 1666464484
transform 1 0 48024 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1666464484
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1666464484
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1666464484
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1666464484
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_560
timestamp 1666464484
transform 1 0 52624 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_572
timestamp 1666464484
transform 1 0 53728 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_584
timestamp 1666464484
transform 1 0 54832 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_596
timestamp 1666464484
transform 1 0 55936 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_603
timestamp 1666464484
transform 1 0 56580 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_615
timestamp 1666464484
transform 1 0 57684 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_623
timestamp 1666464484
transform 1 0 58420 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_22
timestamp 1666464484
transform 1 0 3128 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_34
timestamp 1666464484
transform 1 0 4232 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_46
timestamp 1666464484
transform 1 0 5336 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_58
timestamp 1666464484
transform 1 0 6440 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_89
timestamp 1666464484
transform 1 0 9292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_101
timestamp 1666464484
transform 1 0 10396 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_108
timestamp 1666464484
transform 1 0 11040 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_120
timestamp 1666464484
transform 1 0 12144 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_132
timestamp 1666464484
transform 1 0 13248 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_144
timestamp 1666464484
transform 1 0 14352 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_151
timestamp 1666464484
transform 1 0 14996 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_163
timestamp 1666464484
transform 1 0 16100 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_175
timestamp 1666464484
transform 1 0 17204 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_187
timestamp 1666464484
transform 1 0 18308 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_194
timestamp 1666464484
transform 1 0 18952 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_206
timestamp 1666464484
transform 1 0 20056 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_218
timestamp 1666464484
transform 1 0 21160 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_230
timestamp 1666464484
transform 1 0 22264 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_237
timestamp 1666464484
transform 1 0 22908 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_249
timestamp 1666464484
transform 1 0 24012 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_261
timestamp 1666464484
transform 1 0 25116 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_273
timestamp 1666464484
transform 1 0 26220 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_280
timestamp 1666464484
transform 1 0 26864 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_292
timestamp 1666464484
transform 1 0 27968 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_304
timestamp 1666464484
transform 1 0 29072 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_316
timestamp 1666464484
transform 1 0 30176 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_323
timestamp 1666464484
transform 1 0 30820 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_335
timestamp 1666464484
transform 1 0 31924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_347
timestamp 1666464484
transform 1 0 33028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_359
timestamp 1666464484
transform 1 0 34132 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_366
timestamp 1666464484
transform 1 0 34776 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_378
timestamp 1666464484
transform 1 0 35880 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_390
timestamp 1666464484
transform 1 0 36984 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_402
timestamp 1666464484
transform 1 0 38088 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_409
timestamp 1666464484
transform 1 0 38732 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1666464484
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1666464484
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_445
timestamp 1666464484
transform 1 0 42044 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_452
timestamp 1666464484
transform 1 0 42688 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_464
timestamp 1666464484
transform 1 0 43792 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_476
timestamp 1666464484
transform 1 0 44896 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_488
timestamp 1666464484
transform 1 0 46000 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_495
timestamp 1666464484
transform 1 0 46644 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_507
timestamp 1666464484
transform 1 0 47748 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_519
timestamp 1666464484
transform 1 0 48852 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_531
timestamp 1666464484
transform 1 0 49956 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_538
timestamp 1666464484
transform 1 0 50600 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_550
timestamp 1666464484
transform 1 0 51704 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_562
timestamp 1666464484
transform 1 0 52808 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_574
timestamp 1666464484
transform 1 0 53912 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_581
timestamp 1666464484
transform 1 0 54556 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_593
timestamp 1666464484
transform 1 0 55660 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_605
timestamp 1666464484
transform 1 0 56764 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_617
timestamp 1666464484
transform 1 0 57868 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_624
timestamp 1666464484
transform 1 0 58512 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_44
timestamp 1666464484
transform 1 0 5152 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_56
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_68
timestamp 1666464484
transform 1 0 7360 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_80
timestamp 1666464484
transform 1 0 8464 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_87
timestamp 1666464484
transform 1 0 9108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_99
timestamp 1666464484
transform 1 0 10212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_123
timestamp 1666464484
transform 1 0 12420 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_130
timestamp 1666464484
transform 1 0 13064 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_142
timestamp 1666464484
transform 1 0 14168 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_154
timestamp 1666464484
transform 1 0 15272 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_166
timestamp 1666464484
transform 1 0 16376 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_173
timestamp 1666464484
transform 1 0 17020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_185
timestamp 1666464484
transform 1 0 18124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_197
timestamp 1666464484
transform 1 0 19228 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_209
timestamp 1666464484
transform 1 0 20332 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_216
timestamp 1666464484
transform 1 0 20976 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_228
timestamp 1666464484
transform 1 0 22080 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_240
timestamp 1666464484
transform 1 0 23184 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_252
timestamp 1666464484
transform 1 0 24288 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_259
timestamp 1666464484
transform 1 0 24932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_271
timestamp 1666464484
transform 1 0 26036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_283
timestamp 1666464484
transform 1 0 27140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_295
timestamp 1666464484
transform 1 0 28244 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_302
timestamp 1666464484
transform 1 0 28888 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_314
timestamp 1666464484
transform 1 0 29992 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_326
timestamp 1666464484
transform 1 0 31096 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_338
timestamp 1666464484
transform 1 0 32200 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_345
timestamp 1666464484
transform 1 0 32844 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_357
timestamp 1666464484
transform 1 0 33948 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_369
timestamp 1666464484
transform 1 0 35052 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_381
timestamp 1666464484
transform 1 0 36156 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_388
timestamp 1666464484
transform 1 0 36800 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_400
timestamp 1666464484
transform 1 0 37904 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_412
timestamp 1666464484
transform 1 0 39008 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_424
timestamp 1666464484
transform 1 0 40112 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_431
timestamp 1666464484
transform 1 0 40756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_443
timestamp 1666464484
transform 1 0 41860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_455
timestamp 1666464484
transform 1 0 42964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_467
timestamp 1666464484
transform 1 0 44068 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_474
timestamp 1666464484
transform 1 0 44712 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_486
timestamp 1666464484
transform 1 0 45816 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_498
timestamp 1666464484
transform 1 0 46920 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_510
timestamp 1666464484
transform 1 0 48024 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1666464484
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1666464484
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1666464484
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1666464484
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_560
timestamp 1666464484
transform 1 0 52624 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_572
timestamp 1666464484
transform 1 0 53728 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_584
timestamp 1666464484
transform 1 0 54832 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_596
timestamp 1666464484
transform 1 0 55936 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_603
timestamp 1666464484
transform 1 0 56580 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_615
timestamp 1666464484
transform 1 0 57684 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_623
timestamp 1666464484
transform 1 0 58420 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_15
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_22
timestamp 1666464484
transform 1 0 3128 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_34
timestamp 1666464484
transform 1 0 4232 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_46
timestamp 1666464484
transform 1 0 5336 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_58
timestamp 1666464484
transform 1 0 6440 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_89
timestamp 1666464484
transform 1 0 9292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_101
timestamp 1666464484
transform 1 0 10396 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_108
timestamp 1666464484
transform 1 0 11040 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_120
timestamp 1666464484
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_132
timestamp 1666464484
transform 1 0 13248 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_144
timestamp 1666464484
transform 1 0 14352 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_151
timestamp 1666464484
transform 1 0 14996 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_163
timestamp 1666464484
transform 1 0 16100 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_175
timestamp 1666464484
transform 1 0 17204 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_187
timestamp 1666464484
transform 1 0 18308 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_194
timestamp 1666464484
transform 1 0 18952 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_206
timestamp 1666464484
transform 1 0 20056 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_218
timestamp 1666464484
transform 1 0 21160 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_230
timestamp 1666464484
transform 1 0 22264 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_237
timestamp 1666464484
transform 1 0 22908 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_249
timestamp 1666464484
transform 1 0 24012 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_261
timestamp 1666464484
transform 1 0 25116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_273
timestamp 1666464484
transform 1 0 26220 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_280
timestamp 1666464484
transform 1 0 26864 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_292
timestamp 1666464484
transform 1 0 27968 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_304
timestamp 1666464484
transform 1 0 29072 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_316
timestamp 1666464484
transform 1 0 30176 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_323
timestamp 1666464484
transform 1 0 30820 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_335
timestamp 1666464484
transform 1 0 31924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_347
timestamp 1666464484
transform 1 0 33028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_359
timestamp 1666464484
transform 1 0 34132 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_366
timestamp 1666464484
transform 1 0 34776 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_378
timestamp 1666464484
transform 1 0 35880 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_390
timestamp 1666464484
transform 1 0 36984 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_402
timestamp 1666464484
transform 1 0 38088 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_409
timestamp 1666464484
transform 1 0 38732 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1666464484
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1666464484
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_445
timestamp 1666464484
transform 1 0 42044 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_452
timestamp 1666464484
transform 1 0 42688 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_464
timestamp 1666464484
transform 1 0 43792 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_476
timestamp 1666464484
transform 1 0 44896 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_488
timestamp 1666464484
transform 1 0 46000 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_495
timestamp 1666464484
transform 1 0 46644 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_507
timestamp 1666464484
transform 1 0 47748 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_519
timestamp 1666464484
transform 1 0 48852 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_531
timestamp 1666464484
transform 1 0 49956 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_538
timestamp 1666464484
transform 1 0 50600 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_550
timestamp 1666464484
transform 1 0 51704 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_562
timestamp 1666464484
transform 1 0 52808 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_574
timestamp 1666464484
transform 1 0 53912 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_581
timestamp 1666464484
transform 1 0 54556 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_593
timestamp 1666464484
transform 1 0 55660 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_605
timestamp 1666464484
transform 1 0 56764 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_617
timestamp 1666464484
transform 1 0 57868 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_624
timestamp 1666464484
transform 1 0 58512 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_39
timestamp 1666464484
transform 1 0 4692 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_44
timestamp 1666464484
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_56
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_68
timestamp 1666464484
transform 1 0 7360 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_80
timestamp 1666464484
transform 1 0 8464 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_87
timestamp 1666464484
transform 1 0 9108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_99
timestamp 1666464484
transform 1 0 10212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_123
timestamp 1666464484
transform 1 0 12420 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_130
timestamp 1666464484
transform 1 0 13064 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_142
timestamp 1666464484
transform 1 0 14168 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_154
timestamp 1666464484
transform 1 0 15272 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_166
timestamp 1666464484
transform 1 0 16376 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_173
timestamp 1666464484
transform 1 0 17020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_185
timestamp 1666464484
transform 1 0 18124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_197
timestamp 1666464484
transform 1 0 19228 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_209
timestamp 1666464484
transform 1 0 20332 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_216
timestamp 1666464484
transform 1 0 20976 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_228
timestamp 1666464484
transform 1 0 22080 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_240
timestamp 1666464484
transform 1 0 23184 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_252
timestamp 1666464484
transform 1 0 24288 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_259
timestamp 1666464484
transform 1 0 24932 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_271
timestamp 1666464484
transform 1 0 26036 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_283
timestamp 1666464484
transform 1 0 27140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_295
timestamp 1666464484
transform 1 0 28244 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_302
timestamp 1666464484
transform 1 0 28888 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_314
timestamp 1666464484
transform 1 0 29992 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_326
timestamp 1666464484
transform 1 0 31096 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_338
timestamp 1666464484
transform 1 0 32200 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_345
timestamp 1666464484
transform 1 0 32844 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_357
timestamp 1666464484
transform 1 0 33948 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_369
timestamp 1666464484
transform 1 0 35052 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_381
timestamp 1666464484
transform 1 0 36156 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_388
timestamp 1666464484
transform 1 0 36800 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_400
timestamp 1666464484
transform 1 0 37904 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_412
timestamp 1666464484
transform 1 0 39008 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_424
timestamp 1666464484
transform 1 0 40112 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_431
timestamp 1666464484
transform 1 0 40756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_443
timestamp 1666464484
transform 1 0 41860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_455
timestamp 1666464484
transform 1 0 42964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_467
timestamp 1666464484
transform 1 0 44068 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_474
timestamp 1666464484
transform 1 0 44712 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_486
timestamp 1666464484
transform 1 0 45816 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_498
timestamp 1666464484
transform 1 0 46920 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_510
timestamp 1666464484
transform 1 0 48024 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1666464484
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1666464484
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1666464484
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1666464484
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_560
timestamp 1666464484
transform 1 0 52624 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_572
timestamp 1666464484
transform 1 0 53728 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_584
timestamp 1666464484
transform 1 0 54832 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_596
timestamp 1666464484
transform 1 0 55936 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_603
timestamp 1666464484
transform 1 0 56580 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_615
timestamp 1666464484
transform 1 0 57684 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_623
timestamp 1666464484
transform 1 0 58420 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_22
timestamp 1666464484
transform 1 0 3128 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_34
timestamp 1666464484
transform 1 0 4232 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_46
timestamp 1666464484
transform 1 0 5336 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_58
timestamp 1666464484
transform 1 0 6440 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_89
timestamp 1666464484
transform 1 0 9292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_101
timestamp 1666464484
transform 1 0 10396 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_108
timestamp 1666464484
transform 1 0 11040 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_120
timestamp 1666464484
transform 1 0 12144 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_132
timestamp 1666464484
transform 1 0 13248 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_144
timestamp 1666464484
transform 1 0 14352 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_151
timestamp 1666464484
transform 1 0 14996 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_163
timestamp 1666464484
transform 1 0 16100 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_175
timestamp 1666464484
transform 1 0 17204 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_187
timestamp 1666464484
transform 1 0 18308 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_194
timestamp 1666464484
transform 1 0 18952 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_206
timestamp 1666464484
transform 1 0 20056 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_218
timestamp 1666464484
transform 1 0 21160 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_230
timestamp 1666464484
transform 1 0 22264 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_237
timestamp 1666464484
transform 1 0 22908 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_249
timestamp 1666464484
transform 1 0 24012 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_261
timestamp 1666464484
transform 1 0 25116 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_273
timestamp 1666464484
transform 1 0 26220 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_280
timestamp 1666464484
transform 1 0 26864 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_292
timestamp 1666464484
transform 1 0 27968 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_304
timestamp 1666464484
transform 1 0 29072 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_316
timestamp 1666464484
transform 1 0 30176 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_323
timestamp 1666464484
transform 1 0 30820 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_335
timestamp 1666464484
transform 1 0 31924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_347
timestamp 1666464484
transform 1 0 33028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_359
timestamp 1666464484
transform 1 0 34132 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_366
timestamp 1666464484
transform 1 0 34776 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_378
timestamp 1666464484
transform 1 0 35880 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_390
timestamp 1666464484
transform 1 0 36984 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_402
timestamp 1666464484
transform 1 0 38088 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_409
timestamp 1666464484
transform 1 0 38732 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1666464484
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1666464484
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_445
timestamp 1666464484
transform 1 0 42044 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_452
timestamp 1666464484
transform 1 0 42688 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_464
timestamp 1666464484
transform 1 0 43792 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_476
timestamp 1666464484
transform 1 0 44896 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_488
timestamp 1666464484
transform 1 0 46000 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_495
timestamp 1666464484
transform 1 0 46644 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_507
timestamp 1666464484
transform 1 0 47748 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_519
timestamp 1666464484
transform 1 0 48852 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_531
timestamp 1666464484
transform 1 0 49956 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_538
timestamp 1666464484
transform 1 0 50600 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_550
timestamp 1666464484
transform 1 0 51704 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_562
timestamp 1666464484
transform 1 0 52808 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_574
timestamp 1666464484
transform 1 0 53912 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_581
timestamp 1666464484
transform 1 0 54556 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_593
timestamp 1666464484
transform 1 0 55660 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_605
timestamp 1666464484
transform 1 0 56764 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_617
timestamp 1666464484
transform 1 0 57868 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_624
timestamp 1666464484
transform 1 0 58512 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_39
timestamp 1666464484
transform 1 0 4692 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_44
timestamp 1666464484
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_56
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_68
timestamp 1666464484
transform 1 0 7360 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_80
timestamp 1666464484
transform 1 0 8464 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_87
timestamp 1666464484
transform 1 0 9108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_99
timestamp 1666464484
transform 1 0 10212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_123
timestamp 1666464484
transform 1 0 12420 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_130
timestamp 1666464484
transform 1 0 13064 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_142
timestamp 1666464484
transform 1 0 14168 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_154
timestamp 1666464484
transform 1 0 15272 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_166
timestamp 1666464484
transform 1 0 16376 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_173
timestamp 1666464484
transform 1 0 17020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_185
timestamp 1666464484
transform 1 0 18124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_197
timestamp 1666464484
transform 1 0 19228 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_209
timestamp 1666464484
transform 1 0 20332 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_216
timestamp 1666464484
transform 1 0 20976 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_228
timestamp 1666464484
transform 1 0 22080 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_240
timestamp 1666464484
transform 1 0 23184 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_252
timestamp 1666464484
transform 1 0 24288 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_259
timestamp 1666464484
transform 1 0 24932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_271
timestamp 1666464484
transform 1 0 26036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_283
timestamp 1666464484
transform 1 0 27140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_295
timestamp 1666464484
transform 1 0 28244 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_302
timestamp 1666464484
transform 1 0 28888 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_314
timestamp 1666464484
transform 1 0 29992 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_326
timestamp 1666464484
transform 1 0 31096 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_338
timestamp 1666464484
transform 1 0 32200 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_345
timestamp 1666464484
transform 1 0 32844 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_357
timestamp 1666464484
transform 1 0 33948 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_369
timestamp 1666464484
transform 1 0 35052 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_381
timestamp 1666464484
transform 1 0 36156 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_388
timestamp 1666464484
transform 1 0 36800 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_400
timestamp 1666464484
transform 1 0 37904 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_412
timestamp 1666464484
transform 1 0 39008 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_424
timestamp 1666464484
transform 1 0 40112 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_431
timestamp 1666464484
transform 1 0 40756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_443
timestamp 1666464484
transform 1 0 41860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_455
timestamp 1666464484
transform 1 0 42964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_467
timestamp 1666464484
transform 1 0 44068 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_474
timestamp 1666464484
transform 1 0 44712 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_486
timestamp 1666464484
transform 1 0 45816 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_498
timestamp 1666464484
transform 1 0 46920 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_510
timestamp 1666464484
transform 1 0 48024 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1666464484
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1666464484
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1666464484
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1666464484
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_560
timestamp 1666464484
transform 1 0 52624 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_572
timestamp 1666464484
transform 1 0 53728 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_584
timestamp 1666464484
transform 1 0 54832 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_596
timestamp 1666464484
transform 1 0 55936 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_603
timestamp 1666464484
transform 1 0 56580 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_615
timestamp 1666464484
transform 1 0 57684 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_623
timestamp 1666464484
transform 1 0 58420 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_22
timestamp 1666464484
transform 1 0 3128 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_34
timestamp 1666464484
transform 1 0 4232 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_46
timestamp 1666464484
transform 1 0 5336 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_58
timestamp 1666464484
transform 1 0 6440 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_89
timestamp 1666464484
transform 1 0 9292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_101
timestamp 1666464484
transform 1 0 10396 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_108
timestamp 1666464484
transform 1 0 11040 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_120
timestamp 1666464484
transform 1 0 12144 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_132
timestamp 1666464484
transform 1 0 13248 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_144
timestamp 1666464484
transform 1 0 14352 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_151
timestamp 1666464484
transform 1 0 14996 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_163
timestamp 1666464484
transform 1 0 16100 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_175
timestamp 1666464484
transform 1 0 17204 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_187
timestamp 1666464484
transform 1 0 18308 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_194
timestamp 1666464484
transform 1 0 18952 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_206
timestamp 1666464484
transform 1 0 20056 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_218
timestamp 1666464484
transform 1 0 21160 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_230
timestamp 1666464484
transform 1 0 22264 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_237
timestamp 1666464484
transform 1 0 22908 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_249
timestamp 1666464484
transform 1 0 24012 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_261
timestamp 1666464484
transform 1 0 25116 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_273
timestamp 1666464484
transform 1 0 26220 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_280
timestamp 1666464484
transform 1 0 26864 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_292
timestamp 1666464484
transform 1 0 27968 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_304
timestamp 1666464484
transform 1 0 29072 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_316
timestamp 1666464484
transform 1 0 30176 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_323
timestamp 1666464484
transform 1 0 30820 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_335
timestamp 1666464484
transform 1 0 31924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_347
timestamp 1666464484
transform 1 0 33028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_359
timestamp 1666464484
transform 1 0 34132 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_366
timestamp 1666464484
transform 1 0 34776 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_378
timestamp 1666464484
transform 1 0 35880 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_390
timestamp 1666464484
transform 1 0 36984 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_402
timestamp 1666464484
transform 1 0 38088 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_409
timestamp 1666464484
transform 1 0 38732 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1666464484
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1666464484
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_445
timestamp 1666464484
transform 1 0 42044 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_452
timestamp 1666464484
transform 1 0 42688 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_464
timestamp 1666464484
transform 1 0 43792 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_476
timestamp 1666464484
transform 1 0 44896 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_488
timestamp 1666464484
transform 1 0 46000 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_495
timestamp 1666464484
transform 1 0 46644 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_507
timestamp 1666464484
transform 1 0 47748 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_519
timestamp 1666464484
transform 1 0 48852 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_531
timestamp 1666464484
transform 1 0 49956 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_538
timestamp 1666464484
transform 1 0 50600 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_550
timestamp 1666464484
transform 1 0 51704 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_562
timestamp 1666464484
transform 1 0 52808 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_574
timestamp 1666464484
transform 1 0 53912 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_581
timestamp 1666464484
transform 1 0 54556 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_593
timestamp 1666464484
transform 1 0 55660 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_605
timestamp 1666464484
transform 1 0 56764 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_617
timestamp 1666464484
transform 1 0 57868 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_624
timestamp 1666464484
transform 1 0 58512 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666464484
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1666464484
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_39
timestamp 1666464484
transform 1 0 4692 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_44
timestamp 1666464484
transform 1 0 5152 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_56
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_68
timestamp 1666464484
transform 1 0 7360 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_80
timestamp 1666464484
transform 1 0 8464 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_87
timestamp 1666464484
transform 1 0 9108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_99
timestamp 1666464484
transform 1 0 10212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_123
timestamp 1666464484
transform 1 0 12420 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_130
timestamp 1666464484
transform 1 0 13064 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_142
timestamp 1666464484
transform 1 0 14168 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_154
timestamp 1666464484
transform 1 0 15272 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_166
timestamp 1666464484
transform 1 0 16376 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_173
timestamp 1666464484
transform 1 0 17020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_185
timestamp 1666464484
transform 1 0 18124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_197
timestamp 1666464484
transform 1 0 19228 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_209
timestamp 1666464484
transform 1 0 20332 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_216
timestamp 1666464484
transform 1 0 20976 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_228
timestamp 1666464484
transform 1 0 22080 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_240
timestamp 1666464484
transform 1 0 23184 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_252
timestamp 1666464484
transform 1 0 24288 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_259
timestamp 1666464484
transform 1 0 24932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_271
timestamp 1666464484
transform 1 0 26036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_283
timestamp 1666464484
transform 1 0 27140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_295
timestamp 1666464484
transform 1 0 28244 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_302
timestamp 1666464484
transform 1 0 28888 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_314
timestamp 1666464484
transform 1 0 29992 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_326
timestamp 1666464484
transform 1 0 31096 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_338
timestamp 1666464484
transform 1 0 32200 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_345
timestamp 1666464484
transform 1 0 32844 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_357
timestamp 1666464484
transform 1 0 33948 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_369
timestamp 1666464484
transform 1 0 35052 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_381
timestamp 1666464484
transform 1 0 36156 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_388
timestamp 1666464484
transform 1 0 36800 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_400
timestamp 1666464484
transform 1 0 37904 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_412
timestamp 1666464484
transform 1 0 39008 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_424
timestamp 1666464484
transform 1 0 40112 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_431
timestamp 1666464484
transform 1 0 40756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_443
timestamp 1666464484
transform 1 0 41860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_455
timestamp 1666464484
transform 1 0 42964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_467
timestamp 1666464484
transform 1 0 44068 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_474
timestamp 1666464484
transform 1 0 44712 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_486
timestamp 1666464484
transform 1 0 45816 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_498
timestamp 1666464484
transform 1 0 46920 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_510
timestamp 1666464484
transform 1 0 48024 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1666464484
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1666464484
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1666464484
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1666464484
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_560
timestamp 1666464484
transform 1 0 52624 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_572
timestamp 1666464484
transform 1 0 53728 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_584
timestamp 1666464484
transform 1 0 54832 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_596
timestamp 1666464484
transform 1 0 55936 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_603
timestamp 1666464484
transform 1 0 56580 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_615
timestamp 1666464484
transform 1 0 57684 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_623
timestamp 1666464484
transform 1 0 58420 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_22
timestamp 1666464484
transform 1 0 3128 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_34
timestamp 1666464484
transform 1 0 4232 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_46
timestamp 1666464484
transform 1 0 5336 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_58
timestamp 1666464484
transform 1 0 6440 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_89
timestamp 1666464484
transform 1 0 9292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_101
timestamp 1666464484
transform 1 0 10396 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_108
timestamp 1666464484
transform 1 0 11040 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_120
timestamp 1666464484
transform 1 0 12144 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_132
timestamp 1666464484
transform 1 0 13248 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_144
timestamp 1666464484
transform 1 0 14352 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_151
timestamp 1666464484
transform 1 0 14996 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_163
timestamp 1666464484
transform 1 0 16100 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_175
timestamp 1666464484
transform 1 0 17204 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_187
timestamp 1666464484
transform 1 0 18308 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_194
timestamp 1666464484
transform 1 0 18952 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_206
timestamp 1666464484
transform 1 0 20056 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_218
timestamp 1666464484
transform 1 0 21160 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_230
timestamp 1666464484
transform 1 0 22264 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_237
timestamp 1666464484
transform 1 0 22908 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_249
timestamp 1666464484
transform 1 0 24012 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_261
timestamp 1666464484
transform 1 0 25116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_273
timestamp 1666464484
transform 1 0 26220 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_280
timestamp 1666464484
transform 1 0 26864 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_292
timestamp 1666464484
transform 1 0 27968 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_304
timestamp 1666464484
transform 1 0 29072 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_316
timestamp 1666464484
transform 1 0 30176 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_323
timestamp 1666464484
transform 1 0 30820 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_335
timestamp 1666464484
transform 1 0 31924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_347
timestamp 1666464484
transform 1 0 33028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_359
timestamp 1666464484
transform 1 0 34132 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_366
timestamp 1666464484
transform 1 0 34776 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_378
timestamp 1666464484
transform 1 0 35880 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_390
timestamp 1666464484
transform 1 0 36984 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_402
timestamp 1666464484
transform 1 0 38088 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_409
timestamp 1666464484
transform 1 0 38732 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1666464484
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1666464484
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_445
timestamp 1666464484
transform 1 0 42044 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_452
timestamp 1666464484
transform 1 0 42688 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_464
timestamp 1666464484
transform 1 0 43792 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_476
timestamp 1666464484
transform 1 0 44896 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_488
timestamp 1666464484
transform 1 0 46000 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_495
timestamp 1666464484
transform 1 0 46644 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_507
timestamp 1666464484
transform 1 0 47748 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_519
timestamp 1666464484
transform 1 0 48852 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_531
timestamp 1666464484
transform 1 0 49956 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_538
timestamp 1666464484
transform 1 0 50600 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_550
timestamp 1666464484
transform 1 0 51704 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_562
timestamp 1666464484
transform 1 0 52808 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_574
timestamp 1666464484
transform 1 0 53912 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_581
timestamp 1666464484
transform 1 0 54556 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_593
timestamp 1666464484
transform 1 0 55660 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_605
timestamp 1666464484
transform 1 0 56764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_617
timestamp 1666464484
transform 1 0 57868 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_624
timestamp 1666464484
transform 1 0 58512 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666464484
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666464484
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_39
timestamp 1666464484
transform 1 0 4692 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_44
timestamp 1666464484
transform 1 0 5152 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_56
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_68
timestamp 1666464484
transform 1 0 7360 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_80
timestamp 1666464484
transform 1 0 8464 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_87
timestamp 1666464484
transform 1 0 9108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_99
timestamp 1666464484
transform 1 0 10212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_123
timestamp 1666464484
transform 1 0 12420 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_130
timestamp 1666464484
transform 1 0 13064 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_142
timestamp 1666464484
transform 1 0 14168 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_154
timestamp 1666464484
transform 1 0 15272 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_166
timestamp 1666464484
transform 1 0 16376 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_173
timestamp 1666464484
transform 1 0 17020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_185
timestamp 1666464484
transform 1 0 18124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_197
timestamp 1666464484
transform 1 0 19228 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_209
timestamp 1666464484
transform 1 0 20332 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_216
timestamp 1666464484
transform 1 0 20976 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_228
timestamp 1666464484
transform 1 0 22080 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_240
timestamp 1666464484
transform 1 0 23184 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_252
timestamp 1666464484
transform 1 0 24288 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_259
timestamp 1666464484
transform 1 0 24932 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_271
timestamp 1666464484
transform 1 0 26036 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_283
timestamp 1666464484
transform 1 0 27140 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_295
timestamp 1666464484
transform 1 0 28244 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_302
timestamp 1666464484
transform 1 0 28888 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_314
timestamp 1666464484
transform 1 0 29992 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_326
timestamp 1666464484
transform 1 0 31096 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_338
timestamp 1666464484
transform 1 0 32200 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_345
timestamp 1666464484
transform 1 0 32844 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_357
timestamp 1666464484
transform 1 0 33948 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_369
timestamp 1666464484
transform 1 0 35052 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_381
timestamp 1666464484
transform 1 0 36156 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_388
timestamp 1666464484
transform 1 0 36800 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_400
timestamp 1666464484
transform 1 0 37904 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_412
timestamp 1666464484
transform 1 0 39008 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_424
timestamp 1666464484
transform 1 0 40112 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_431
timestamp 1666464484
transform 1 0 40756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_443
timestamp 1666464484
transform 1 0 41860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_455
timestamp 1666464484
transform 1 0 42964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_467
timestamp 1666464484
transform 1 0 44068 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_474
timestamp 1666464484
transform 1 0 44712 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_486
timestamp 1666464484
transform 1 0 45816 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_498
timestamp 1666464484
transform 1 0 46920 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_510
timestamp 1666464484
transform 1 0 48024 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1666464484
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1666464484
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1666464484
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1666464484
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_560
timestamp 1666464484
transform 1 0 52624 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_572
timestamp 1666464484
transform 1 0 53728 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_584
timestamp 1666464484
transform 1 0 54832 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_596
timestamp 1666464484
transform 1 0 55936 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_603
timestamp 1666464484
transform 1 0 56580 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_615
timestamp 1666464484
transform 1 0 57684 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_623
timestamp 1666464484
transform 1 0 58420 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_15
timestamp 1666464484
transform 1 0 2484 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_22
timestamp 1666464484
transform 1 0 3128 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_34
timestamp 1666464484
transform 1 0 4232 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_46
timestamp 1666464484
transform 1 0 5336 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_58
timestamp 1666464484
transform 1 0 6440 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_89
timestamp 1666464484
transform 1 0 9292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_101
timestamp 1666464484
transform 1 0 10396 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_108
timestamp 1666464484
transform 1 0 11040 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_120
timestamp 1666464484
transform 1 0 12144 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_132
timestamp 1666464484
transform 1 0 13248 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_144
timestamp 1666464484
transform 1 0 14352 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_151
timestamp 1666464484
transform 1 0 14996 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_163
timestamp 1666464484
transform 1 0 16100 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_175
timestamp 1666464484
transform 1 0 17204 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_187
timestamp 1666464484
transform 1 0 18308 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_194
timestamp 1666464484
transform 1 0 18952 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_206
timestamp 1666464484
transform 1 0 20056 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_218
timestamp 1666464484
transform 1 0 21160 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_230
timestamp 1666464484
transform 1 0 22264 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_237
timestamp 1666464484
transform 1 0 22908 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_249
timestamp 1666464484
transform 1 0 24012 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_261
timestamp 1666464484
transform 1 0 25116 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_273
timestamp 1666464484
transform 1 0 26220 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_280
timestamp 1666464484
transform 1 0 26864 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_292
timestamp 1666464484
transform 1 0 27968 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_304
timestamp 1666464484
transform 1 0 29072 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_316
timestamp 1666464484
transform 1 0 30176 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_323
timestamp 1666464484
transform 1 0 30820 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_335
timestamp 1666464484
transform 1 0 31924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_347
timestamp 1666464484
transform 1 0 33028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_359
timestamp 1666464484
transform 1 0 34132 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_366
timestamp 1666464484
transform 1 0 34776 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_378
timestamp 1666464484
transform 1 0 35880 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_390
timestamp 1666464484
transform 1 0 36984 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_402
timestamp 1666464484
transform 1 0 38088 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_409
timestamp 1666464484
transform 1 0 38732 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1666464484
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1666464484
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_445
timestamp 1666464484
transform 1 0 42044 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_452
timestamp 1666464484
transform 1 0 42688 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_464
timestamp 1666464484
transform 1 0 43792 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_476
timestamp 1666464484
transform 1 0 44896 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_488
timestamp 1666464484
transform 1 0 46000 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_495
timestamp 1666464484
transform 1 0 46644 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_507
timestamp 1666464484
transform 1 0 47748 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_519
timestamp 1666464484
transform 1 0 48852 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_531
timestamp 1666464484
transform 1 0 49956 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_538
timestamp 1666464484
transform 1 0 50600 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_550
timestamp 1666464484
transform 1 0 51704 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_562
timestamp 1666464484
transform 1 0 52808 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_574
timestamp 1666464484
transform 1 0 53912 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_581
timestamp 1666464484
transform 1 0 54556 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_593
timestamp 1666464484
transform 1 0 55660 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_605
timestamp 1666464484
transform 1 0 56764 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_617
timestamp 1666464484
transform 1 0 57868 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_624
timestamp 1666464484
transform 1 0 58512 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_44
timestamp 1666464484
transform 1 0 5152 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_56
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_68
timestamp 1666464484
transform 1 0 7360 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_80
timestamp 1666464484
transform 1 0 8464 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_87
timestamp 1666464484
transform 1 0 9108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_99
timestamp 1666464484
transform 1 0 10212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_123
timestamp 1666464484
transform 1 0 12420 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_130
timestamp 1666464484
transform 1 0 13064 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_142
timestamp 1666464484
transform 1 0 14168 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_154
timestamp 1666464484
transform 1 0 15272 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_166
timestamp 1666464484
transform 1 0 16376 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_173
timestamp 1666464484
transform 1 0 17020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_185
timestamp 1666464484
transform 1 0 18124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_197
timestamp 1666464484
transform 1 0 19228 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_209
timestamp 1666464484
transform 1 0 20332 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_216
timestamp 1666464484
transform 1 0 20976 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_228
timestamp 1666464484
transform 1 0 22080 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_240
timestamp 1666464484
transform 1 0 23184 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_252
timestamp 1666464484
transform 1 0 24288 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_259
timestamp 1666464484
transform 1 0 24932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_271
timestamp 1666464484
transform 1 0 26036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_283
timestamp 1666464484
transform 1 0 27140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_295
timestamp 1666464484
transform 1 0 28244 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_302
timestamp 1666464484
transform 1 0 28888 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_314
timestamp 1666464484
transform 1 0 29992 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_326
timestamp 1666464484
transform 1 0 31096 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_338
timestamp 1666464484
transform 1 0 32200 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_345
timestamp 1666464484
transform 1 0 32844 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_357
timestamp 1666464484
transform 1 0 33948 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_369
timestamp 1666464484
transform 1 0 35052 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_381
timestamp 1666464484
transform 1 0 36156 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_388
timestamp 1666464484
transform 1 0 36800 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_400
timestamp 1666464484
transform 1 0 37904 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_412
timestamp 1666464484
transform 1 0 39008 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_424
timestamp 1666464484
transform 1 0 40112 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_431
timestamp 1666464484
transform 1 0 40756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_443
timestamp 1666464484
transform 1 0 41860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_455
timestamp 1666464484
transform 1 0 42964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_467
timestamp 1666464484
transform 1 0 44068 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_474
timestamp 1666464484
transform 1 0 44712 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_486
timestamp 1666464484
transform 1 0 45816 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_498
timestamp 1666464484
transform 1 0 46920 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_510
timestamp 1666464484
transform 1 0 48024 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1666464484
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1666464484
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1666464484
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1666464484
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_560
timestamp 1666464484
transform 1 0 52624 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_572
timestamp 1666464484
transform 1 0 53728 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_584
timestamp 1666464484
transform 1 0 54832 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_596
timestamp 1666464484
transform 1 0 55936 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_603
timestamp 1666464484
transform 1 0 56580 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_615
timestamp 1666464484
transform 1 0 57684 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_623
timestamp 1666464484
transform 1 0 58420 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_22
timestamp 1666464484
transform 1 0 3128 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_34
timestamp 1666464484
transform 1 0 4232 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_46
timestamp 1666464484
transform 1 0 5336 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_58
timestamp 1666464484
transform 1 0 6440 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_77
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_89
timestamp 1666464484
transform 1 0 9292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_101
timestamp 1666464484
transform 1 0 10396 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_108
timestamp 1666464484
transform 1 0 11040 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_120
timestamp 1666464484
transform 1 0 12144 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_132
timestamp 1666464484
transform 1 0 13248 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_144
timestamp 1666464484
transform 1 0 14352 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_151
timestamp 1666464484
transform 1 0 14996 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_163
timestamp 1666464484
transform 1 0 16100 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_175
timestamp 1666464484
transform 1 0 17204 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_187
timestamp 1666464484
transform 1 0 18308 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_194
timestamp 1666464484
transform 1 0 18952 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_206
timestamp 1666464484
transform 1 0 20056 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_218
timestamp 1666464484
transform 1 0 21160 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_230
timestamp 1666464484
transform 1 0 22264 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_237
timestamp 1666464484
transform 1 0 22908 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_249
timestamp 1666464484
transform 1 0 24012 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_261
timestamp 1666464484
transform 1 0 25116 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_273
timestamp 1666464484
transform 1 0 26220 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_280
timestamp 1666464484
transform 1 0 26864 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_292
timestamp 1666464484
transform 1 0 27968 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_304
timestamp 1666464484
transform 1 0 29072 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_316
timestamp 1666464484
transform 1 0 30176 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_323
timestamp 1666464484
transform 1 0 30820 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_335
timestamp 1666464484
transform 1 0 31924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_347
timestamp 1666464484
transform 1 0 33028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_359
timestamp 1666464484
transform 1 0 34132 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_366
timestamp 1666464484
transform 1 0 34776 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_378
timestamp 1666464484
transform 1 0 35880 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_390
timestamp 1666464484
transform 1 0 36984 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_402
timestamp 1666464484
transform 1 0 38088 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_409
timestamp 1666464484
transform 1 0 38732 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1666464484
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1666464484
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_445
timestamp 1666464484
transform 1 0 42044 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_452
timestamp 1666464484
transform 1 0 42688 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_464
timestamp 1666464484
transform 1 0 43792 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_476
timestamp 1666464484
transform 1 0 44896 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_488
timestamp 1666464484
transform 1 0 46000 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_495
timestamp 1666464484
transform 1 0 46644 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_507
timestamp 1666464484
transform 1 0 47748 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_519
timestamp 1666464484
transform 1 0 48852 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_531
timestamp 1666464484
transform 1 0 49956 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_538
timestamp 1666464484
transform 1 0 50600 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_550
timestamp 1666464484
transform 1 0 51704 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_562
timestamp 1666464484
transform 1 0 52808 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_574
timestamp 1666464484
transform 1 0 53912 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_581
timestamp 1666464484
transform 1 0 54556 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_593
timestamp 1666464484
transform 1 0 55660 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_605
timestamp 1666464484
transform 1 0 56764 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_617
timestamp 1666464484
transform 1 0 57868 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_624
timestamp 1666464484
transform 1 0 58512 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666464484
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666464484
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_39
timestamp 1666464484
transform 1 0 4692 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_44
timestamp 1666464484
transform 1 0 5152 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_56
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_68
timestamp 1666464484
transform 1 0 7360 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_80
timestamp 1666464484
transform 1 0 8464 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_87
timestamp 1666464484
transform 1 0 9108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_99
timestamp 1666464484
transform 1 0 10212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_123
timestamp 1666464484
transform 1 0 12420 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_130
timestamp 1666464484
transform 1 0 13064 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_142
timestamp 1666464484
transform 1 0 14168 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_154
timestamp 1666464484
transform 1 0 15272 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_166
timestamp 1666464484
transform 1 0 16376 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_173
timestamp 1666464484
transform 1 0 17020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_185
timestamp 1666464484
transform 1 0 18124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_197
timestamp 1666464484
transform 1 0 19228 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_209
timestamp 1666464484
transform 1 0 20332 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_216
timestamp 1666464484
transform 1 0 20976 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_228
timestamp 1666464484
transform 1 0 22080 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_240
timestamp 1666464484
transform 1 0 23184 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_252
timestamp 1666464484
transform 1 0 24288 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_259
timestamp 1666464484
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_271
timestamp 1666464484
transform 1 0 26036 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_283
timestamp 1666464484
transform 1 0 27140 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_295
timestamp 1666464484
transform 1 0 28244 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_302
timestamp 1666464484
transform 1 0 28888 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_314
timestamp 1666464484
transform 1 0 29992 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_326
timestamp 1666464484
transform 1 0 31096 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_338
timestamp 1666464484
transform 1 0 32200 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_345
timestamp 1666464484
transform 1 0 32844 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_357
timestamp 1666464484
transform 1 0 33948 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_369
timestamp 1666464484
transform 1 0 35052 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_381
timestamp 1666464484
transform 1 0 36156 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_388
timestamp 1666464484
transform 1 0 36800 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_400
timestamp 1666464484
transform 1 0 37904 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_412
timestamp 1666464484
transform 1 0 39008 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_424
timestamp 1666464484
transform 1 0 40112 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_431
timestamp 1666464484
transform 1 0 40756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_443
timestamp 1666464484
transform 1 0 41860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_455
timestamp 1666464484
transform 1 0 42964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_467
timestamp 1666464484
transform 1 0 44068 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_474
timestamp 1666464484
transform 1 0 44712 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_486
timestamp 1666464484
transform 1 0 45816 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_498
timestamp 1666464484
transform 1 0 46920 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_510
timestamp 1666464484
transform 1 0 48024 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1666464484
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1666464484
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1666464484
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1666464484
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_560
timestamp 1666464484
transform 1 0 52624 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_572
timestamp 1666464484
transform 1 0 53728 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_584
timestamp 1666464484
transform 1 0 54832 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_596
timestamp 1666464484
transform 1 0 55936 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_603
timestamp 1666464484
transform 1 0 56580 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_615
timestamp 1666464484
transform 1 0 57684 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_623
timestamp 1666464484
transform 1 0 58420 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_15
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_22
timestamp 1666464484
transform 1 0 3128 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_34
timestamp 1666464484
transform 1 0 4232 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_46
timestamp 1666464484
transform 1 0 5336 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_58
timestamp 1666464484
transform 1 0 6440 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_89
timestamp 1666464484
transform 1 0 9292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_101
timestamp 1666464484
transform 1 0 10396 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_108
timestamp 1666464484
transform 1 0 11040 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_120
timestamp 1666464484
transform 1 0 12144 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_132
timestamp 1666464484
transform 1 0 13248 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_144
timestamp 1666464484
transform 1 0 14352 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_151
timestamp 1666464484
transform 1 0 14996 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_163
timestamp 1666464484
transform 1 0 16100 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_175
timestamp 1666464484
transform 1 0 17204 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_187
timestamp 1666464484
transform 1 0 18308 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_194
timestamp 1666464484
transform 1 0 18952 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_206
timestamp 1666464484
transform 1 0 20056 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_218
timestamp 1666464484
transform 1 0 21160 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_230
timestamp 1666464484
transform 1 0 22264 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_237
timestamp 1666464484
transform 1 0 22908 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_249
timestamp 1666464484
transform 1 0 24012 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_261
timestamp 1666464484
transform 1 0 25116 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_273
timestamp 1666464484
transform 1 0 26220 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_280
timestamp 1666464484
transform 1 0 26864 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_292
timestamp 1666464484
transform 1 0 27968 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_304
timestamp 1666464484
transform 1 0 29072 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_316
timestamp 1666464484
transform 1 0 30176 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_323
timestamp 1666464484
transform 1 0 30820 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_335
timestamp 1666464484
transform 1 0 31924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_347
timestamp 1666464484
transform 1 0 33028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_359
timestamp 1666464484
transform 1 0 34132 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_366
timestamp 1666464484
transform 1 0 34776 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_378
timestamp 1666464484
transform 1 0 35880 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_390
timestamp 1666464484
transform 1 0 36984 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_402
timestamp 1666464484
transform 1 0 38088 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_409
timestamp 1666464484
transform 1 0 38732 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1666464484
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1666464484
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_445
timestamp 1666464484
transform 1 0 42044 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_452
timestamp 1666464484
transform 1 0 42688 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_464
timestamp 1666464484
transform 1 0 43792 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_476
timestamp 1666464484
transform 1 0 44896 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_488
timestamp 1666464484
transform 1 0 46000 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_495
timestamp 1666464484
transform 1 0 46644 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_507
timestamp 1666464484
transform 1 0 47748 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_519
timestamp 1666464484
transform 1 0 48852 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_531
timestamp 1666464484
transform 1 0 49956 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_538
timestamp 1666464484
transform 1 0 50600 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_550
timestamp 1666464484
transform 1 0 51704 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_562
timestamp 1666464484
transform 1 0 52808 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_574
timestamp 1666464484
transform 1 0 53912 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_581
timestamp 1666464484
transform 1 0 54556 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_593
timestamp 1666464484
transform 1 0 55660 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_605
timestamp 1666464484
transform 1 0 56764 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_617
timestamp 1666464484
transform 1 0 57868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_624
timestamp 1666464484
transform 1 0 58512 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_44
timestamp 1666464484
transform 1 0 5152 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_56
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_68
timestamp 1666464484
transform 1 0 7360 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_80
timestamp 1666464484
transform 1 0 8464 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_87
timestamp 1666464484
transform 1 0 9108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_99
timestamp 1666464484
transform 1 0 10212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_111
timestamp 1666464484
transform 1 0 11316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_123
timestamp 1666464484
transform 1 0 12420 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_130
timestamp 1666464484
transform 1 0 13064 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_142
timestamp 1666464484
transform 1 0 14168 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_154
timestamp 1666464484
transform 1 0 15272 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_166
timestamp 1666464484
transform 1 0 16376 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_173
timestamp 1666464484
transform 1 0 17020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_185
timestamp 1666464484
transform 1 0 18124 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_197
timestamp 1666464484
transform 1 0 19228 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_209
timestamp 1666464484
transform 1 0 20332 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_216
timestamp 1666464484
transform 1 0 20976 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_228
timestamp 1666464484
transform 1 0 22080 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_240
timestamp 1666464484
transform 1 0 23184 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_252
timestamp 1666464484
transform 1 0 24288 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_259
timestamp 1666464484
transform 1 0 24932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_271
timestamp 1666464484
transform 1 0 26036 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_283
timestamp 1666464484
transform 1 0 27140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_295
timestamp 1666464484
transform 1 0 28244 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_302
timestamp 1666464484
transform 1 0 28888 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_314
timestamp 1666464484
transform 1 0 29992 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_326
timestamp 1666464484
transform 1 0 31096 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_338
timestamp 1666464484
transform 1 0 32200 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_345
timestamp 1666464484
transform 1 0 32844 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_357
timestamp 1666464484
transform 1 0 33948 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_369
timestamp 1666464484
transform 1 0 35052 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_381
timestamp 1666464484
transform 1 0 36156 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_388
timestamp 1666464484
transform 1 0 36800 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_400
timestamp 1666464484
transform 1 0 37904 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_412
timestamp 1666464484
transform 1 0 39008 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_424
timestamp 1666464484
transform 1 0 40112 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_431
timestamp 1666464484
transform 1 0 40756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_443
timestamp 1666464484
transform 1 0 41860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_455
timestamp 1666464484
transform 1 0 42964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_467
timestamp 1666464484
transform 1 0 44068 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_474
timestamp 1666464484
transform 1 0 44712 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_486
timestamp 1666464484
transform 1 0 45816 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_498
timestamp 1666464484
transform 1 0 46920 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_510
timestamp 1666464484
transform 1 0 48024 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1666464484
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1666464484
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1666464484
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1666464484
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_560
timestamp 1666464484
transform 1 0 52624 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_572
timestamp 1666464484
transform 1 0 53728 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_584
timestamp 1666464484
transform 1 0 54832 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_596
timestamp 1666464484
transform 1 0 55936 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_603
timestamp 1666464484
transform 1 0 56580 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_615
timestamp 1666464484
transform 1 0 57684 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_623
timestamp 1666464484
transform 1 0 58420 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_22
timestamp 1666464484
transform 1 0 3128 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_34
timestamp 1666464484
transform 1 0 4232 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_46
timestamp 1666464484
transform 1 0 5336 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_58
timestamp 1666464484
transform 1 0 6440 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666464484
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_77
timestamp 1666464484
transform 1 0 8188 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_89
timestamp 1666464484
transform 1 0 9292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_101
timestamp 1666464484
transform 1 0 10396 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_108
timestamp 1666464484
transform 1 0 11040 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_120
timestamp 1666464484
transform 1 0 12144 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_132
timestamp 1666464484
transform 1 0 13248 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_144
timestamp 1666464484
transform 1 0 14352 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_151
timestamp 1666464484
transform 1 0 14996 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_163
timestamp 1666464484
transform 1 0 16100 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_175
timestamp 1666464484
transform 1 0 17204 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_187
timestamp 1666464484
transform 1 0 18308 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_194
timestamp 1666464484
transform 1 0 18952 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_206
timestamp 1666464484
transform 1 0 20056 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_218
timestamp 1666464484
transform 1 0 21160 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_230
timestamp 1666464484
transform 1 0 22264 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_237
timestamp 1666464484
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_249
timestamp 1666464484
transform 1 0 24012 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_261
timestamp 1666464484
transform 1 0 25116 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_273
timestamp 1666464484
transform 1 0 26220 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_280
timestamp 1666464484
transform 1 0 26864 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_292
timestamp 1666464484
transform 1 0 27968 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_304
timestamp 1666464484
transform 1 0 29072 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_316
timestamp 1666464484
transform 1 0 30176 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_323
timestamp 1666464484
transform 1 0 30820 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_335
timestamp 1666464484
transform 1 0 31924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_347
timestamp 1666464484
transform 1 0 33028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_359
timestamp 1666464484
transform 1 0 34132 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_366
timestamp 1666464484
transform 1 0 34776 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_378
timestamp 1666464484
transform 1 0 35880 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_390
timestamp 1666464484
transform 1 0 36984 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_402
timestamp 1666464484
transform 1 0 38088 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_409
timestamp 1666464484
transform 1 0 38732 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1666464484
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1666464484
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_445
timestamp 1666464484
transform 1 0 42044 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_452
timestamp 1666464484
transform 1 0 42688 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_464
timestamp 1666464484
transform 1 0 43792 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_476
timestamp 1666464484
transform 1 0 44896 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_488
timestamp 1666464484
transform 1 0 46000 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_495
timestamp 1666464484
transform 1 0 46644 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_507
timestamp 1666464484
transform 1 0 47748 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_519
timestamp 1666464484
transform 1 0 48852 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_531
timestamp 1666464484
transform 1 0 49956 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_538
timestamp 1666464484
transform 1 0 50600 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_550
timestamp 1666464484
transform 1 0 51704 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_562
timestamp 1666464484
transform 1 0 52808 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_574
timestamp 1666464484
transform 1 0 53912 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_581
timestamp 1666464484
transform 1 0 54556 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_593
timestamp 1666464484
transform 1 0 55660 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_605
timestamp 1666464484
transform 1 0 56764 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_617
timestamp 1666464484
transform 1 0 57868 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_624
timestamp 1666464484
transform 1 0 58512 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_39
timestamp 1666464484
transform 1 0 4692 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1666464484
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_56
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_68
timestamp 1666464484
transform 1 0 7360 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_80
timestamp 1666464484
transform 1 0 8464 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_87
timestamp 1666464484
transform 1 0 9108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_99
timestamp 1666464484
transform 1 0 10212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_111
timestamp 1666464484
transform 1 0 11316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_123
timestamp 1666464484
transform 1 0 12420 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_130
timestamp 1666464484
transform 1 0 13064 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_142
timestamp 1666464484
transform 1 0 14168 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_154
timestamp 1666464484
transform 1 0 15272 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_166
timestamp 1666464484
transform 1 0 16376 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_173
timestamp 1666464484
transform 1 0 17020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_185
timestamp 1666464484
transform 1 0 18124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_197
timestamp 1666464484
transform 1 0 19228 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_209
timestamp 1666464484
transform 1 0 20332 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_216
timestamp 1666464484
transform 1 0 20976 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_228
timestamp 1666464484
transform 1 0 22080 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_240
timestamp 1666464484
transform 1 0 23184 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_252
timestamp 1666464484
transform 1 0 24288 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_259
timestamp 1666464484
transform 1 0 24932 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_271
timestamp 1666464484
transform 1 0 26036 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_283
timestamp 1666464484
transform 1 0 27140 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_295
timestamp 1666464484
transform 1 0 28244 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_302
timestamp 1666464484
transform 1 0 28888 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_314
timestamp 1666464484
transform 1 0 29992 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_326
timestamp 1666464484
transform 1 0 31096 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_338
timestamp 1666464484
transform 1 0 32200 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_345
timestamp 1666464484
transform 1 0 32844 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_357
timestamp 1666464484
transform 1 0 33948 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_369
timestamp 1666464484
transform 1 0 35052 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_381
timestamp 1666464484
transform 1 0 36156 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_388
timestamp 1666464484
transform 1 0 36800 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_400
timestamp 1666464484
transform 1 0 37904 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_412
timestamp 1666464484
transform 1 0 39008 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_424
timestamp 1666464484
transform 1 0 40112 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_431
timestamp 1666464484
transform 1 0 40756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_443
timestamp 1666464484
transform 1 0 41860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_455
timestamp 1666464484
transform 1 0 42964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_467
timestamp 1666464484
transform 1 0 44068 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_474
timestamp 1666464484
transform 1 0 44712 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_486
timestamp 1666464484
transform 1 0 45816 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_498
timestamp 1666464484
transform 1 0 46920 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_510
timestamp 1666464484
transform 1 0 48024 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1666464484
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1666464484
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1666464484
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1666464484
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_560
timestamp 1666464484
transform 1 0 52624 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_572
timestamp 1666464484
transform 1 0 53728 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_584
timestamp 1666464484
transform 1 0 54832 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_596
timestamp 1666464484
transform 1 0 55936 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_603
timestamp 1666464484
transform 1 0 56580 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_615
timestamp 1666464484
transform 1 0 57684 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_623
timestamp 1666464484
transform 1 0 58420 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_15
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_22
timestamp 1666464484
transform 1 0 3128 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_34
timestamp 1666464484
transform 1 0 4232 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_46
timestamp 1666464484
transform 1 0 5336 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_58
timestamp 1666464484
transform 1 0 6440 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_77
timestamp 1666464484
transform 1 0 8188 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_89
timestamp 1666464484
transform 1 0 9292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_101
timestamp 1666464484
transform 1 0 10396 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_108
timestamp 1666464484
transform 1 0 11040 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_120
timestamp 1666464484
transform 1 0 12144 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_132
timestamp 1666464484
transform 1 0 13248 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_144
timestamp 1666464484
transform 1 0 14352 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_151
timestamp 1666464484
transform 1 0 14996 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_163
timestamp 1666464484
transform 1 0 16100 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_175
timestamp 1666464484
transform 1 0 17204 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_187
timestamp 1666464484
transform 1 0 18308 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_194
timestamp 1666464484
transform 1 0 18952 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_206
timestamp 1666464484
transform 1 0 20056 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_218
timestamp 1666464484
transform 1 0 21160 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_230
timestamp 1666464484
transform 1 0 22264 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_237
timestamp 1666464484
transform 1 0 22908 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_249
timestamp 1666464484
transform 1 0 24012 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_261
timestamp 1666464484
transform 1 0 25116 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_273
timestamp 1666464484
transform 1 0 26220 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_280
timestamp 1666464484
transform 1 0 26864 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_292
timestamp 1666464484
transform 1 0 27968 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_304
timestamp 1666464484
transform 1 0 29072 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_316
timestamp 1666464484
transform 1 0 30176 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_323
timestamp 1666464484
transform 1 0 30820 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_335
timestamp 1666464484
transform 1 0 31924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_347
timestamp 1666464484
transform 1 0 33028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_359
timestamp 1666464484
transform 1 0 34132 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_366
timestamp 1666464484
transform 1 0 34776 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_378
timestamp 1666464484
transform 1 0 35880 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_390
timestamp 1666464484
transform 1 0 36984 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_402
timestamp 1666464484
transform 1 0 38088 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_409
timestamp 1666464484
transform 1 0 38732 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1666464484
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1666464484
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_445
timestamp 1666464484
transform 1 0 42044 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_452
timestamp 1666464484
transform 1 0 42688 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_464
timestamp 1666464484
transform 1 0 43792 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_476
timestamp 1666464484
transform 1 0 44896 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_488
timestamp 1666464484
transform 1 0 46000 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_495
timestamp 1666464484
transform 1 0 46644 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_507
timestamp 1666464484
transform 1 0 47748 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_519
timestamp 1666464484
transform 1 0 48852 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_531
timestamp 1666464484
transform 1 0 49956 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_538
timestamp 1666464484
transform 1 0 50600 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_550
timestamp 1666464484
transform 1 0 51704 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_562
timestamp 1666464484
transform 1 0 52808 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_574
timestamp 1666464484
transform 1 0 53912 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_581
timestamp 1666464484
transform 1 0 54556 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_593
timestamp 1666464484
transform 1 0 55660 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_605
timestamp 1666464484
transform 1 0 56764 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_617
timestamp 1666464484
transform 1 0 57868 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_624
timestamp 1666464484
transform 1 0 58512 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_44
timestamp 1666464484
transform 1 0 5152 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_56
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_68
timestamp 1666464484
transform 1 0 7360 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_80
timestamp 1666464484
transform 1 0 8464 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_87
timestamp 1666464484
transform 1 0 9108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_99
timestamp 1666464484
transform 1 0 10212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_111
timestamp 1666464484
transform 1 0 11316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_123
timestamp 1666464484
transform 1 0 12420 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_130
timestamp 1666464484
transform 1 0 13064 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_142
timestamp 1666464484
transform 1 0 14168 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_154
timestamp 1666464484
transform 1 0 15272 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_166
timestamp 1666464484
transform 1 0 16376 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_173
timestamp 1666464484
transform 1 0 17020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_185
timestamp 1666464484
transform 1 0 18124 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_197
timestamp 1666464484
transform 1 0 19228 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_209
timestamp 1666464484
transform 1 0 20332 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_216
timestamp 1666464484
transform 1 0 20976 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_228
timestamp 1666464484
transform 1 0 22080 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_240
timestamp 1666464484
transform 1 0 23184 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_252
timestamp 1666464484
transform 1 0 24288 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_259
timestamp 1666464484
transform 1 0 24932 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_271
timestamp 1666464484
transform 1 0 26036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_283
timestamp 1666464484
transform 1 0 27140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_295
timestamp 1666464484
transform 1 0 28244 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_302
timestamp 1666464484
transform 1 0 28888 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_314
timestamp 1666464484
transform 1 0 29992 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_326
timestamp 1666464484
transform 1 0 31096 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_338
timestamp 1666464484
transform 1 0 32200 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_345
timestamp 1666464484
transform 1 0 32844 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_357
timestamp 1666464484
transform 1 0 33948 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_369
timestamp 1666464484
transform 1 0 35052 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_381
timestamp 1666464484
transform 1 0 36156 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_388
timestamp 1666464484
transform 1 0 36800 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_400
timestamp 1666464484
transform 1 0 37904 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_412
timestamp 1666464484
transform 1 0 39008 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_424
timestamp 1666464484
transform 1 0 40112 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_431
timestamp 1666464484
transform 1 0 40756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_443
timestamp 1666464484
transform 1 0 41860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_455
timestamp 1666464484
transform 1 0 42964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_467
timestamp 1666464484
transform 1 0 44068 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_474
timestamp 1666464484
transform 1 0 44712 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_486
timestamp 1666464484
transform 1 0 45816 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_498
timestamp 1666464484
transform 1 0 46920 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_510
timestamp 1666464484
transform 1 0 48024 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1666464484
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1666464484
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1666464484
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1666464484
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_560
timestamp 1666464484
transform 1 0 52624 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_572
timestamp 1666464484
transform 1 0 53728 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_584
timestamp 1666464484
transform 1 0 54832 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_596
timestamp 1666464484
transform 1 0 55936 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_603
timestamp 1666464484
transform 1 0 56580 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_615
timestamp 1666464484
transform 1 0 57684 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_623
timestamp 1666464484
transform 1 0 58420 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_15
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_22
timestamp 1666464484
transform 1 0 3128 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_34
timestamp 1666464484
transform 1 0 4232 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_46
timestamp 1666464484
transform 1 0 5336 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_58
timestamp 1666464484
transform 1 0 6440 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_89
timestamp 1666464484
transform 1 0 9292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_101
timestamp 1666464484
transform 1 0 10396 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_108
timestamp 1666464484
transform 1 0 11040 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_120
timestamp 1666464484
transform 1 0 12144 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_132
timestamp 1666464484
transform 1 0 13248 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_144
timestamp 1666464484
transform 1 0 14352 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_151
timestamp 1666464484
transform 1 0 14996 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_163
timestamp 1666464484
transform 1 0 16100 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_175
timestamp 1666464484
transform 1 0 17204 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_187
timestamp 1666464484
transform 1 0 18308 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_194
timestamp 1666464484
transform 1 0 18952 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_206
timestamp 1666464484
transform 1 0 20056 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_218
timestamp 1666464484
transform 1 0 21160 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_230
timestamp 1666464484
transform 1 0 22264 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_237
timestamp 1666464484
transform 1 0 22908 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_249
timestamp 1666464484
transform 1 0 24012 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_261
timestamp 1666464484
transform 1 0 25116 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_273
timestamp 1666464484
transform 1 0 26220 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_280
timestamp 1666464484
transform 1 0 26864 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_292
timestamp 1666464484
transform 1 0 27968 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_304
timestamp 1666464484
transform 1 0 29072 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_316
timestamp 1666464484
transform 1 0 30176 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_323
timestamp 1666464484
transform 1 0 30820 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_335
timestamp 1666464484
transform 1 0 31924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_347
timestamp 1666464484
transform 1 0 33028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_359
timestamp 1666464484
transform 1 0 34132 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_366
timestamp 1666464484
transform 1 0 34776 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_378
timestamp 1666464484
transform 1 0 35880 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_390
timestamp 1666464484
transform 1 0 36984 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_402
timestamp 1666464484
transform 1 0 38088 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_409
timestamp 1666464484
transform 1 0 38732 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1666464484
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1666464484
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_445
timestamp 1666464484
transform 1 0 42044 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_452
timestamp 1666464484
transform 1 0 42688 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_464
timestamp 1666464484
transform 1 0 43792 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_476
timestamp 1666464484
transform 1 0 44896 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_488
timestamp 1666464484
transform 1 0 46000 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_495
timestamp 1666464484
transform 1 0 46644 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_507
timestamp 1666464484
transform 1 0 47748 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_519
timestamp 1666464484
transform 1 0 48852 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_531
timestamp 1666464484
transform 1 0 49956 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_538
timestamp 1666464484
transform 1 0 50600 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_550
timestamp 1666464484
transform 1 0 51704 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_562
timestamp 1666464484
transform 1 0 52808 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_574
timestamp 1666464484
transform 1 0 53912 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_581
timestamp 1666464484
transform 1 0 54556 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_593
timestamp 1666464484
transform 1 0 55660 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_605
timestamp 1666464484
transform 1 0 56764 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_617
timestamp 1666464484
transform 1 0 57868 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_624
timestamp 1666464484
transform 1 0 58512 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_44
timestamp 1666464484
transform 1 0 5152 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_56
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_68
timestamp 1666464484
transform 1 0 7360 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_80
timestamp 1666464484
transform 1 0 8464 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_87
timestamp 1666464484
transform 1 0 9108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_99
timestamp 1666464484
transform 1 0 10212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_123
timestamp 1666464484
transform 1 0 12420 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_130
timestamp 1666464484
transform 1 0 13064 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_142
timestamp 1666464484
transform 1 0 14168 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_154
timestamp 1666464484
transform 1 0 15272 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_166
timestamp 1666464484
transform 1 0 16376 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_173
timestamp 1666464484
transform 1 0 17020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_185
timestamp 1666464484
transform 1 0 18124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_197
timestamp 1666464484
transform 1 0 19228 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_209
timestamp 1666464484
transform 1 0 20332 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_216
timestamp 1666464484
transform 1 0 20976 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_228
timestamp 1666464484
transform 1 0 22080 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_240
timestamp 1666464484
transform 1 0 23184 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_252
timestamp 1666464484
transform 1 0 24288 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_259
timestamp 1666464484
transform 1 0 24932 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_271
timestamp 1666464484
transform 1 0 26036 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_283
timestamp 1666464484
transform 1 0 27140 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_295
timestamp 1666464484
transform 1 0 28244 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_302
timestamp 1666464484
transform 1 0 28888 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_314
timestamp 1666464484
transform 1 0 29992 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_326
timestamp 1666464484
transform 1 0 31096 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_338
timestamp 1666464484
transform 1 0 32200 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_345
timestamp 1666464484
transform 1 0 32844 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_357
timestamp 1666464484
transform 1 0 33948 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_369
timestamp 1666464484
transform 1 0 35052 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_381
timestamp 1666464484
transform 1 0 36156 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_388
timestamp 1666464484
transform 1 0 36800 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_400
timestamp 1666464484
transform 1 0 37904 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_412
timestamp 1666464484
transform 1 0 39008 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_424
timestamp 1666464484
transform 1 0 40112 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_431
timestamp 1666464484
transform 1 0 40756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_443
timestamp 1666464484
transform 1 0 41860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_455
timestamp 1666464484
transform 1 0 42964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_467
timestamp 1666464484
transform 1 0 44068 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_474
timestamp 1666464484
transform 1 0 44712 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_486
timestamp 1666464484
transform 1 0 45816 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_498
timestamp 1666464484
transform 1 0 46920 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_510
timestamp 1666464484
transform 1 0 48024 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1666464484
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1666464484
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1666464484
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1666464484
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_560
timestamp 1666464484
transform 1 0 52624 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_572
timestamp 1666464484
transform 1 0 53728 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_584
timestamp 1666464484
transform 1 0 54832 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_596
timestamp 1666464484
transform 1 0 55936 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_603
timestamp 1666464484
transform 1 0 56580 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_615
timestamp 1666464484
transform 1 0 57684 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_623
timestamp 1666464484
transform 1 0 58420 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_15
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_22
timestamp 1666464484
transform 1 0 3128 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_34
timestamp 1666464484
transform 1 0 4232 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_46
timestamp 1666464484
transform 1 0 5336 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_58
timestamp 1666464484
transform 1 0 6440 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_89
timestamp 1666464484
transform 1 0 9292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_101
timestamp 1666464484
transform 1 0 10396 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_108
timestamp 1666464484
transform 1 0 11040 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_120
timestamp 1666464484
transform 1 0 12144 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_132
timestamp 1666464484
transform 1 0 13248 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_144
timestamp 1666464484
transform 1 0 14352 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_151
timestamp 1666464484
transform 1 0 14996 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_163
timestamp 1666464484
transform 1 0 16100 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_175
timestamp 1666464484
transform 1 0 17204 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_187
timestamp 1666464484
transform 1 0 18308 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_194
timestamp 1666464484
transform 1 0 18952 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_206
timestamp 1666464484
transform 1 0 20056 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_218
timestamp 1666464484
transform 1 0 21160 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_230
timestamp 1666464484
transform 1 0 22264 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_237
timestamp 1666464484
transform 1 0 22908 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_249
timestamp 1666464484
transform 1 0 24012 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_261
timestamp 1666464484
transform 1 0 25116 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_273
timestamp 1666464484
transform 1 0 26220 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_280
timestamp 1666464484
transform 1 0 26864 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_292
timestamp 1666464484
transform 1 0 27968 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_304
timestamp 1666464484
transform 1 0 29072 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_316
timestamp 1666464484
transform 1 0 30176 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_323
timestamp 1666464484
transform 1 0 30820 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_335
timestamp 1666464484
transform 1 0 31924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_347
timestamp 1666464484
transform 1 0 33028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_359
timestamp 1666464484
transform 1 0 34132 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_366
timestamp 1666464484
transform 1 0 34776 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_378
timestamp 1666464484
transform 1 0 35880 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_390
timestamp 1666464484
transform 1 0 36984 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_402
timestamp 1666464484
transform 1 0 38088 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_409
timestamp 1666464484
transform 1 0 38732 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1666464484
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1666464484
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_445
timestamp 1666464484
transform 1 0 42044 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_452
timestamp 1666464484
transform 1 0 42688 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_464
timestamp 1666464484
transform 1 0 43792 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_476
timestamp 1666464484
transform 1 0 44896 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_488
timestamp 1666464484
transform 1 0 46000 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_495
timestamp 1666464484
transform 1 0 46644 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_507
timestamp 1666464484
transform 1 0 47748 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_519
timestamp 1666464484
transform 1 0 48852 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_531
timestamp 1666464484
transform 1 0 49956 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_538
timestamp 1666464484
transform 1 0 50600 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_550
timestamp 1666464484
transform 1 0 51704 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_562
timestamp 1666464484
transform 1 0 52808 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_574
timestamp 1666464484
transform 1 0 53912 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_581
timestamp 1666464484
transform 1 0 54556 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_593
timestamp 1666464484
transform 1 0 55660 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_605
timestamp 1666464484
transform 1 0 56764 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_617
timestamp 1666464484
transform 1 0 57868 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_624
timestamp 1666464484
transform 1 0 58512 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666464484
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666464484
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_39
timestamp 1666464484
transform 1 0 4692 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_44
timestamp 1666464484
transform 1 0 5152 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_56
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_68
timestamp 1666464484
transform 1 0 7360 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_80
timestamp 1666464484
transform 1 0 8464 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_87
timestamp 1666464484
transform 1 0 9108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_99
timestamp 1666464484
transform 1 0 10212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_111
timestamp 1666464484
transform 1 0 11316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_123
timestamp 1666464484
transform 1 0 12420 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_130
timestamp 1666464484
transform 1 0 13064 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_142
timestamp 1666464484
transform 1 0 14168 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_154
timestamp 1666464484
transform 1 0 15272 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_166
timestamp 1666464484
transform 1 0 16376 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_173
timestamp 1666464484
transform 1 0 17020 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_185
timestamp 1666464484
transform 1 0 18124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_197
timestamp 1666464484
transform 1 0 19228 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_209
timestamp 1666464484
transform 1 0 20332 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_216
timestamp 1666464484
transform 1 0 20976 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_228
timestamp 1666464484
transform 1 0 22080 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_240
timestamp 1666464484
transform 1 0 23184 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_252
timestamp 1666464484
transform 1 0 24288 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_259
timestamp 1666464484
transform 1 0 24932 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_271
timestamp 1666464484
transform 1 0 26036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_283
timestamp 1666464484
transform 1 0 27140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_295
timestamp 1666464484
transform 1 0 28244 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_302
timestamp 1666464484
transform 1 0 28888 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_314
timestamp 1666464484
transform 1 0 29992 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_326
timestamp 1666464484
transform 1 0 31096 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_338
timestamp 1666464484
transform 1 0 32200 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_345
timestamp 1666464484
transform 1 0 32844 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_357
timestamp 1666464484
transform 1 0 33948 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_369
timestamp 1666464484
transform 1 0 35052 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_381
timestamp 1666464484
transform 1 0 36156 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_388
timestamp 1666464484
transform 1 0 36800 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_400
timestamp 1666464484
transform 1 0 37904 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_412
timestamp 1666464484
transform 1 0 39008 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_424
timestamp 1666464484
transform 1 0 40112 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_431
timestamp 1666464484
transform 1 0 40756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_443
timestamp 1666464484
transform 1 0 41860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_455
timestamp 1666464484
transform 1 0 42964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_467
timestamp 1666464484
transform 1 0 44068 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_474
timestamp 1666464484
transform 1 0 44712 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_486
timestamp 1666464484
transform 1 0 45816 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_498
timestamp 1666464484
transform 1 0 46920 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_510
timestamp 1666464484
transform 1 0 48024 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1666464484
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1666464484
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1666464484
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1666464484
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_560
timestamp 1666464484
transform 1 0 52624 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_572
timestamp 1666464484
transform 1 0 53728 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_584
timestamp 1666464484
transform 1 0 54832 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_596
timestamp 1666464484
transform 1 0 55936 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_603
timestamp 1666464484
transform 1 0 56580 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_615
timestamp 1666464484
transform 1 0 57684 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_623
timestamp 1666464484
transform 1 0 58420 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_15
timestamp 1666464484
transform 1 0 2484 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_22
timestamp 1666464484
transform 1 0 3128 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_34
timestamp 1666464484
transform 1 0 4232 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_46
timestamp 1666464484
transform 1 0 5336 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_58
timestamp 1666464484
transform 1 0 6440 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_89
timestamp 1666464484
transform 1 0 9292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_101
timestamp 1666464484
transform 1 0 10396 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_108
timestamp 1666464484
transform 1 0 11040 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_120
timestamp 1666464484
transform 1 0 12144 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_132
timestamp 1666464484
transform 1 0 13248 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_144
timestamp 1666464484
transform 1 0 14352 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_151
timestamp 1666464484
transform 1 0 14996 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_163
timestamp 1666464484
transform 1 0 16100 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_175
timestamp 1666464484
transform 1 0 17204 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_187
timestamp 1666464484
transform 1 0 18308 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_194
timestamp 1666464484
transform 1 0 18952 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_206
timestamp 1666464484
transform 1 0 20056 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_218
timestamp 1666464484
transform 1 0 21160 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_230
timestamp 1666464484
transform 1 0 22264 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_237
timestamp 1666464484
transform 1 0 22908 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_249
timestamp 1666464484
transform 1 0 24012 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_261
timestamp 1666464484
transform 1 0 25116 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_273
timestamp 1666464484
transform 1 0 26220 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_280
timestamp 1666464484
transform 1 0 26864 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_292
timestamp 1666464484
transform 1 0 27968 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_304
timestamp 1666464484
transform 1 0 29072 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_316
timestamp 1666464484
transform 1 0 30176 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_323
timestamp 1666464484
transform 1 0 30820 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_335
timestamp 1666464484
transform 1 0 31924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_347
timestamp 1666464484
transform 1 0 33028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_359
timestamp 1666464484
transform 1 0 34132 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_366
timestamp 1666464484
transform 1 0 34776 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_378
timestamp 1666464484
transform 1 0 35880 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_390
timestamp 1666464484
transform 1 0 36984 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_402
timestamp 1666464484
transform 1 0 38088 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_409
timestamp 1666464484
transform 1 0 38732 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1666464484
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1666464484
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_445
timestamp 1666464484
transform 1 0 42044 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_452
timestamp 1666464484
transform 1 0 42688 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_464
timestamp 1666464484
transform 1 0 43792 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_476
timestamp 1666464484
transform 1 0 44896 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_488
timestamp 1666464484
transform 1 0 46000 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_495
timestamp 1666464484
transform 1 0 46644 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_507
timestamp 1666464484
transform 1 0 47748 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_519
timestamp 1666464484
transform 1 0 48852 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_531
timestamp 1666464484
transform 1 0 49956 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_538
timestamp 1666464484
transform 1 0 50600 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_550
timestamp 1666464484
transform 1 0 51704 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_562
timestamp 1666464484
transform 1 0 52808 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_574
timestamp 1666464484
transform 1 0 53912 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_581
timestamp 1666464484
transform 1 0 54556 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_593
timestamp 1666464484
transform 1 0 55660 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_605
timestamp 1666464484
transform 1 0 56764 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_617
timestamp 1666464484
transform 1 0 57868 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_624
timestamp 1666464484
transform 1 0 58512 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_39
timestamp 1666464484
transform 1 0 4692 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_44
timestamp 1666464484
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_56
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_68
timestamp 1666464484
transform 1 0 7360 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_80
timestamp 1666464484
transform 1 0 8464 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_87
timestamp 1666464484
transform 1 0 9108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_99
timestamp 1666464484
transform 1 0 10212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_123
timestamp 1666464484
transform 1 0 12420 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_130
timestamp 1666464484
transform 1 0 13064 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_142
timestamp 1666464484
transform 1 0 14168 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_154
timestamp 1666464484
transform 1 0 15272 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_166
timestamp 1666464484
transform 1 0 16376 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_173
timestamp 1666464484
transform 1 0 17020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_185
timestamp 1666464484
transform 1 0 18124 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_197
timestamp 1666464484
transform 1 0 19228 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_209
timestamp 1666464484
transform 1 0 20332 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_216
timestamp 1666464484
transform 1 0 20976 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_228
timestamp 1666464484
transform 1 0 22080 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_240
timestamp 1666464484
transform 1 0 23184 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_252
timestamp 1666464484
transform 1 0 24288 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_259
timestamp 1666464484
transform 1 0 24932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_271
timestamp 1666464484
transform 1 0 26036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_283
timestamp 1666464484
transform 1 0 27140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_295
timestamp 1666464484
transform 1 0 28244 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_302
timestamp 1666464484
transform 1 0 28888 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_314
timestamp 1666464484
transform 1 0 29992 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_326
timestamp 1666464484
transform 1 0 31096 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_338
timestamp 1666464484
transform 1 0 32200 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_345
timestamp 1666464484
transform 1 0 32844 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_357
timestamp 1666464484
transform 1 0 33948 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_369
timestamp 1666464484
transform 1 0 35052 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_381
timestamp 1666464484
transform 1 0 36156 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_388
timestamp 1666464484
transform 1 0 36800 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_400
timestamp 1666464484
transform 1 0 37904 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_412
timestamp 1666464484
transform 1 0 39008 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_424
timestamp 1666464484
transform 1 0 40112 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_431
timestamp 1666464484
transform 1 0 40756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_443
timestamp 1666464484
transform 1 0 41860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_455
timestamp 1666464484
transform 1 0 42964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_467
timestamp 1666464484
transform 1 0 44068 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_474
timestamp 1666464484
transform 1 0 44712 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_486
timestamp 1666464484
transform 1 0 45816 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_498
timestamp 1666464484
transform 1 0 46920 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_510
timestamp 1666464484
transform 1 0 48024 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1666464484
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1666464484
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1666464484
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1666464484
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_560
timestamp 1666464484
transform 1 0 52624 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_572
timestamp 1666464484
transform 1 0 53728 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_584
timestamp 1666464484
transform 1 0 54832 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_596
timestamp 1666464484
transform 1 0 55936 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_603
timestamp 1666464484
transform 1 0 56580 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_615
timestamp 1666464484
transform 1 0 57684 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_623
timestamp 1666464484
transform 1 0 58420 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_15
timestamp 1666464484
transform 1 0 2484 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_22
timestamp 1666464484
transform 1 0 3128 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_34
timestamp 1666464484
transform 1 0 4232 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_46
timestamp 1666464484
transform 1 0 5336 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_58
timestamp 1666464484
transform 1 0 6440 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666464484
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_89
timestamp 1666464484
transform 1 0 9292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_101
timestamp 1666464484
transform 1 0 10396 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_108
timestamp 1666464484
transform 1 0 11040 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_120
timestamp 1666464484
transform 1 0 12144 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_132
timestamp 1666464484
transform 1 0 13248 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_144
timestamp 1666464484
transform 1 0 14352 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_151
timestamp 1666464484
transform 1 0 14996 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_163
timestamp 1666464484
transform 1 0 16100 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_175
timestamp 1666464484
transform 1 0 17204 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_187
timestamp 1666464484
transform 1 0 18308 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_194
timestamp 1666464484
transform 1 0 18952 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_206
timestamp 1666464484
transform 1 0 20056 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_218
timestamp 1666464484
transform 1 0 21160 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_230
timestamp 1666464484
transform 1 0 22264 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_237
timestamp 1666464484
transform 1 0 22908 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_249
timestamp 1666464484
transform 1 0 24012 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_261
timestamp 1666464484
transform 1 0 25116 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_273
timestamp 1666464484
transform 1 0 26220 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_280
timestamp 1666464484
transform 1 0 26864 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_292
timestamp 1666464484
transform 1 0 27968 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_304
timestamp 1666464484
transform 1 0 29072 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_316
timestamp 1666464484
transform 1 0 30176 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_323
timestamp 1666464484
transform 1 0 30820 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_335
timestamp 1666464484
transform 1 0 31924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_347
timestamp 1666464484
transform 1 0 33028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_359
timestamp 1666464484
transform 1 0 34132 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_366
timestamp 1666464484
transform 1 0 34776 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_378
timestamp 1666464484
transform 1 0 35880 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_390
timestamp 1666464484
transform 1 0 36984 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_402
timestamp 1666464484
transform 1 0 38088 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_409
timestamp 1666464484
transform 1 0 38732 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1666464484
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1666464484
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_445
timestamp 1666464484
transform 1 0 42044 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_452
timestamp 1666464484
transform 1 0 42688 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_464
timestamp 1666464484
transform 1 0 43792 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_476
timestamp 1666464484
transform 1 0 44896 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_488
timestamp 1666464484
transform 1 0 46000 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_495
timestamp 1666464484
transform 1 0 46644 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_507
timestamp 1666464484
transform 1 0 47748 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_519
timestamp 1666464484
transform 1 0 48852 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_531
timestamp 1666464484
transform 1 0 49956 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_538
timestamp 1666464484
transform 1 0 50600 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_550
timestamp 1666464484
transform 1 0 51704 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_562
timestamp 1666464484
transform 1 0 52808 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_574
timestamp 1666464484
transform 1 0 53912 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_581
timestamp 1666464484
transform 1 0 54556 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_593
timestamp 1666464484
transform 1 0 55660 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_605
timestamp 1666464484
transform 1 0 56764 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_617
timestamp 1666464484
transform 1 0 57868 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_624
timestamp 1666464484
transform 1 0 58512 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666464484
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1666464484
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_39
timestamp 1666464484
transform 1 0 4692 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_44
timestamp 1666464484
transform 1 0 5152 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_56
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_68
timestamp 1666464484
transform 1 0 7360 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_80
timestamp 1666464484
transform 1 0 8464 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_87
timestamp 1666464484
transform 1 0 9108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_99
timestamp 1666464484
transform 1 0 10212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_111
timestamp 1666464484
transform 1 0 11316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_123
timestamp 1666464484
transform 1 0 12420 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_130
timestamp 1666464484
transform 1 0 13064 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_142
timestamp 1666464484
transform 1 0 14168 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_154
timestamp 1666464484
transform 1 0 15272 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_166
timestamp 1666464484
transform 1 0 16376 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_173
timestamp 1666464484
transform 1 0 17020 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_185
timestamp 1666464484
transform 1 0 18124 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_197
timestamp 1666464484
transform 1 0 19228 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_209
timestamp 1666464484
transform 1 0 20332 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_216
timestamp 1666464484
transform 1 0 20976 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_228
timestamp 1666464484
transform 1 0 22080 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_240
timestamp 1666464484
transform 1 0 23184 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_252
timestamp 1666464484
transform 1 0 24288 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_259
timestamp 1666464484
transform 1 0 24932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_271
timestamp 1666464484
transform 1 0 26036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_283
timestamp 1666464484
transform 1 0 27140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_295
timestamp 1666464484
transform 1 0 28244 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_302
timestamp 1666464484
transform 1 0 28888 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_314
timestamp 1666464484
transform 1 0 29992 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_326
timestamp 1666464484
transform 1 0 31096 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_338
timestamp 1666464484
transform 1 0 32200 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_345
timestamp 1666464484
transform 1 0 32844 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_357
timestamp 1666464484
transform 1 0 33948 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_369
timestamp 1666464484
transform 1 0 35052 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_381
timestamp 1666464484
transform 1 0 36156 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_388
timestamp 1666464484
transform 1 0 36800 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_400
timestamp 1666464484
transform 1 0 37904 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_412
timestamp 1666464484
transform 1 0 39008 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_424
timestamp 1666464484
transform 1 0 40112 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_431
timestamp 1666464484
transform 1 0 40756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_443
timestamp 1666464484
transform 1 0 41860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_455
timestamp 1666464484
transform 1 0 42964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_467
timestamp 1666464484
transform 1 0 44068 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_474
timestamp 1666464484
transform 1 0 44712 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_486
timestamp 1666464484
transform 1 0 45816 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_498
timestamp 1666464484
transform 1 0 46920 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_510
timestamp 1666464484
transform 1 0 48024 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1666464484
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1666464484
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1666464484
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1666464484
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_560
timestamp 1666464484
transform 1 0 52624 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_572
timestamp 1666464484
transform 1 0 53728 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_584
timestamp 1666464484
transform 1 0 54832 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_596
timestamp 1666464484
transform 1 0 55936 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_603
timestamp 1666464484
transform 1 0 56580 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_615
timestamp 1666464484
transform 1 0 57684 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_623
timestamp 1666464484
transform 1 0 58420 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_15
timestamp 1666464484
transform 1 0 2484 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_22
timestamp 1666464484
transform 1 0 3128 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_34
timestamp 1666464484
transform 1 0 4232 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_46
timestamp 1666464484
transform 1 0 5336 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_58
timestamp 1666464484
transform 1 0 6440 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666464484
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_77
timestamp 1666464484
transform 1 0 8188 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_89
timestamp 1666464484
transform 1 0 9292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_101
timestamp 1666464484
transform 1 0 10396 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_108
timestamp 1666464484
transform 1 0 11040 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_120
timestamp 1666464484
transform 1 0 12144 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_132
timestamp 1666464484
transform 1 0 13248 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_144
timestamp 1666464484
transform 1 0 14352 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_151
timestamp 1666464484
transform 1 0 14996 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_163
timestamp 1666464484
transform 1 0 16100 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_175
timestamp 1666464484
transform 1 0 17204 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_187
timestamp 1666464484
transform 1 0 18308 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_194
timestamp 1666464484
transform 1 0 18952 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_206
timestamp 1666464484
transform 1 0 20056 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_218
timestamp 1666464484
transform 1 0 21160 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_230
timestamp 1666464484
transform 1 0 22264 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_237
timestamp 1666464484
transform 1 0 22908 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_249
timestamp 1666464484
transform 1 0 24012 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_261
timestamp 1666464484
transform 1 0 25116 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_273
timestamp 1666464484
transform 1 0 26220 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_280
timestamp 1666464484
transform 1 0 26864 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_292
timestamp 1666464484
transform 1 0 27968 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_304
timestamp 1666464484
transform 1 0 29072 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_316
timestamp 1666464484
transform 1 0 30176 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_323
timestamp 1666464484
transform 1 0 30820 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_335
timestamp 1666464484
transform 1 0 31924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_347
timestamp 1666464484
transform 1 0 33028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_359
timestamp 1666464484
transform 1 0 34132 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_366
timestamp 1666464484
transform 1 0 34776 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_378
timestamp 1666464484
transform 1 0 35880 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_390
timestamp 1666464484
transform 1 0 36984 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_402
timestamp 1666464484
transform 1 0 38088 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_409
timestamp 1666464484
transform 1 0 38732 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1666464484
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1666464484
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_445
timestamp 1666464484
transform 1 0 42044 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_452
timestamp 1666464484
transform 1 0 42688 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_464
timestamp 1666464484
transform 1 0 43792 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_476
timestamp 1666464484
transform 1 0 44896 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_488
timestamp 1666464484
transform 1 0 46000 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_495
timestamp 1666464484
transform 1 0 46644 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_507
timestamp 1666464484
transform 1 0 47748 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_519
timestamp 1666464484
transform 1 0 48852 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_531
timestamp 1666464484
transform 1 0 49956 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_538
timestamp 1666464484
transform 1 0 50600 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_550
timestamp 1666464484
transform 1 0 51704 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_562
timestamp 1666464484
transform 1 0 52808 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_574
timestamp 1666464484
transform 1 0 53912 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_581
timestamp 1666464484
transform 1 0 54556 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_593
timestamp 1666464484
transform 1 0 55660 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_605
timestamp 1666464484
transform 1 0 56764 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_617
timestamp 1666464484
transform 1 0 57868 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_624
timestamp 1666464484
transform 1 0 58512 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666464484
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666464484
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_39
timestamp 1666464484
transform 1 0 4692 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_44
timestamp 1666464484
transform 1 0 5152 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_56
timestamp 1666464484
transform 1 0 6256 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_68
timestamp 1666464484
transform 1 0 7360 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_80
timestamp 1666464484
transform 1 0 8464 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_87
timestamp 1666464484
transform 1 0 9108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_99
timestamp 1666464484
transform 1 0 10212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_111
timestamp 1666464484
transform 1 0 11316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_123
timestamp 1666464484
transform 1 0 12420 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_130
timestamp 1666464484
transform 1 0 13064 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_142
timestamp 1666464484
transform 1 0 14168 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_154
timestamp 1666464484
transform 1 0 15272 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_166
timestamp 1666464484
transform 1 0 16376 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_173
timestamp 1666464484
transform 1 0 17020 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_185
timestamp 1666464484
transform 1 0 18124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_197
timestamp 1666464484
transform 1 0 19228 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_209
timestamp 1666464484
transform 1 0 20332 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_216
timestamp 1666464484
transform 1 0 20976 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_228
timestamp 1666464484
transform 1 0 22080 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_240
timestamp 1666464484
transform 1 0 23184 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_252
timestamp 1666464484
transform 1 0 24288 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_259
timestamp 1666464484
transform 1 0 24932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_271
timestamp 1666464484
transform 1 0 26036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_283
timestamp 1666464484
transform 1 0 27140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_295
timestamp 1666464484
transform 1 0 28244 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_302
timestamp 1666464484
transform 1 0 28888 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_314
timestamp 1666464484
transform 1 0 29992 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_326
timestamp 1666464484
transform 1 0 31096 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_338
timestamp 1666464484
transform 1 0 32200 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_345
timestamp 1666464484
transform 1 0 32844 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_357
timestamp 1666464484
transform 1 0 33948 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_369
timestamp 1666464484
transform 1 0 35052 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_381
timestamp 1666464484
transform 1 0 36156 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_388
timestamp 1666464484
transform 1 0 36800 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_400
timestamp 1666464484
transform 1 0 37904 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_412
timestamp 1666464484
transform 1 0 39008 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_424
timestamp 1666464484
transform 1 0 40112 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_431
timestamp 1666464484
transform 1 0 40756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_443
timestamp 1666464484
transform 1 0 41860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_455
timestamp 1666464484
transform 1 0 42964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_467
timestamp 1666464484
transform 1 0 44068 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_474
timestamp 1666464484
transform 1 0 44712 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_486
timestamp 1666464484
transform 1 0 45816 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_498
timestamp 1666464484
transform 1 0 46920 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_510
timestamp 1666464484
transform 1 0 48024 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1666464484
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1666464484
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1666464484
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1666464484
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_560
timestamp 1666464484
transform 1 0 52624 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_572
timestamp 1666464484
transform 1 0 53728 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_584
timestamp 1666464484
transform 1 0 54832 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_596
timestamp 1666464484
transform 1 0 55936 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_603
timestamp 1666464484
transform 1 0 56580 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_615
timestamp 1666464484
transform 1 0 57684 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_623
timestamp 1666464484
transform 1 0 58420 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_15
timestamp 1666464484
transform 1 0 2484 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_22
timestamp 1666464484
transform 1 0 3128 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_34
timestamp 1666464484
transform 1 0 4232 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_46
timestamp 1666464484
transform 1 0 5336 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_58
timestamp 1666464484
transform 1 0 6440 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666464484
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_77
timestamp 1666464484
transform 1 0 8188 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_89
timestamp 1666464484
transform 1 0 9292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_101
timestamp 1666464484
transform 1 0 10396 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_108
timestamp 1666464484
transform 1 0 11040 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_120
timestamp 1666464484
transform 1 0 12144 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_132
timestamp 1666464484
transform 1 0 13248 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_144
timestamp 1666464484
transform 1 0 14352 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_151
timestamp 1666464484
transform 1 0 14996 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_163
timestamp 1666464484
transform 1 0 16100 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_175
timestamp 1666464484
transform 1 0 17204 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_187
timestamp 1666464484
transform 1 0 18308 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_194
timestamp 1666464484
transform 1 0 18952 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_206
timestamp 1666464484
transform 1 0 20056 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_218
timestamp 1666464484
transform 1 0 21160 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_230
timestamp 1666464484
transform 1 0 22264 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_237
timestamp 1666464484
transform 1 0 22908 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_249
timestamp 1666464484
transform 1 0 24012 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_261
timestamp 1666464484
transform 1 0 25116 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_273
timestamp 1666464484
transform 1 0 26220 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_280
timestamp 1666464484
transform 1 0 26864 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_292
timestamp 1666464484
transform 1 0 27968 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_304
timestamp 1666464484
transform 1 0 29072 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_316
timestamp 1666464484
transform 1 0 30176 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_323
timestamp 1666464484
transform 1 0 30820 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_335
timestamp 1666464484
transform 1 0 31924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_347
timestamp 1666464484
transform 1 0 33028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_359
timestamp 1666464484
transform 1 0 34132 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_366
timestamp 1666464484
transform 1 0 34776 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_378
timestamp 1666464484
transform 1 0 35880 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_390
timestamp 1666464484
transform 1 0 36984 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_402
timestamp 1666464484
transform 1 0 38088 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_409
timestamp 1666464484
transform 1 0 38732 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1666464484
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1666464484
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_445
timestamp 1666464484
transform 1 0 42044 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_452
timestamp 1666464484
transform 1 0 42688 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_464
timestamp 1666464484
transform 1 0 43792 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_476
timestamp 1666464484
transform 1 0 44896 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_488
timestamp 1666464484
transform 1 0 46000 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_495
timestamp 1666464484
transform 1 0 46644 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_507
timestamp 1666464484
transform 1 0 47748 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_519
timestamp 1666464484
transform 1 0 48852 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_531
timestamp 1666464484
transform 1 0 49956 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_538
timestamp 1666464484
transform 1 0 50600 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_550
timestamp 1666464484
transform 1 0 51704 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_562
timestamp 1666464484
transform 1 0 52808 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_574
timestamp 1666464484
transform 1 0 53912 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_581
timestamp 1666464484
transform 1 0 54556 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_593
timestamp 1666464484
transform 1 0 55660 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_605
timestamp 1666464484
transform 1 0 56764 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_617
timestamp 1666464484
transform 1 0 57868 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_624
timestamp 1666464484
transform 1 0 58512 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666464484
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1666464484
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_39
timestamp 1666464484
transform 1 0 4692 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_44
timestamp 1666464484
transform 1 0 5152 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_56
timestamp 1666464484
transform 1 0 6256 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_68
timestamp 1666464484
transform 1 0 7360 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_80
timestamp 1666464484
transform 1 0 8464 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_87
timestamp 1666464484
transform 1 0 9108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_99
timestamp 1666464484
transform 1 0 10212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_111
timestamp 1666464484
transform 1 0 11316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_123
timestamp 1666464484
transform 1 0 12420 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_130
timestamp 1666464484
transform 1 0 13064 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_142
timestamp 1666464484
transform 1 0 14168 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_154
timestamp 1666464484
transform 1 0 15272 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_166
timestamp 1666464484
transform 1 0 16376 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_173
timestamp 1666464484
transform 1 0 17020 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_185
timestamp 1666464484
transform 1 0 18124 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_197
timestamp 1666464484
transform 1 0 19228 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_209
timestamp 1666464484
transform 1 0 20332 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_216
timestamp 1666464484
transform 1 0 20976 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_228
timestamp 1666464484
transform 1 0 22080 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_240
timestamp 1666464484
transform 1 0 23184 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_252
timestamp 1666464484
transform 1 0 24288 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_259
timestamp 1666464484
transform 1 0 24932 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_271
timestamp 1666464484
transform 1 0 26036 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_283
timestamp 1666464484
transform 1 0 27140 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_295
timestamp 1666464484
transform 1 0 28244 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_302
timestamp 1666464484
transform 1 0 28888 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_314
timestamp 1666464484
transform 1 0 29992 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_326
timestamp 1666464484
transform 1 0 31096 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_338
timestamp 1666464484
transform 1 0 32200 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_345
timestamp 1666464484
transform 1 0 32844 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_357
timestamp 1666464484
transform 1 0 33948 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_369
timestamp 1666464484
transform 1 0 35052 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_381
timestamp 1666464484
transform 1 0 36156 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_388
timestamp 1666464484
transform 1 0 36800 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_400
timestamp 1666464484
transform 1 0 37904 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_412
timestamp 1666464484
transform 1 0 39008 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_424
timestamp 1666464484
transform 1 0 40112 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_431
timestamp 1666464484
transform 1 0 40756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_443
timestamp 1666464484
transform 1 0 41860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_455
timestamp 1666464484
transform 1 0 42964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_467
timestamp 1666464484
transform 1 0 44068 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_474
timestamp 1666464484
transform 1 0 44712 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_486
timestamp 1666464484
transform 1 0 45816 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_498
timestamp 1666464484
transform 1 0 46920 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_510
timestamp 1666464484
transform 1 0 48024 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1666464484
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1666464484
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1666464484
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1666464484
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_560
timestamp 1666464484
transform 1 0 52624 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_572
timestamp 1666464484
transform 1 0 53728 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_584
timestamp 1666464484
transform 1 0 54832 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_596
timestamp 1666464484
transform 1 0 55936 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_603
timestamp 1666464484
transform 1 0 56580 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_615
timestamp 1666464484
transform 1 0 57684 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_623
timestamp 1666464484
transform 1 0 58420 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_15
timestamp 1666464484
transform 1 0 2484 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_22
timestamp 1666464484
transform 1 0 3128 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_34
timestamp 1666464484
transform 1 0 4232 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_46
timestamp 1666464484
transform 1 0 5336 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_58
timestamp 1666464484
transform 1 0 6440 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1666464484
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_77
timestamp 1666464484
transform 1 0 8188 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_89
timestamp 1666464484
transform 1 0 9292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_101
timestamp 1666464484
transform 1 0 10396 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_108
timestamp 1666464484
transform 1 0 11040 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_120
timestamp 1666464484
transform 1 0 12144 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_132
timestamp 1666464484
transform 1 0 13248 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_144
timestamp 1666464484
transform 1 0 14352 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_151
timestamp 1666464484
transform 1 0 14996 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_163
timestamp 1666464484
transform 1 0 16100 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_175
timestamp 1666464484
transform 1 0 17204 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_187
timestamp 1666464484
transform 1 0 18308 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_194
timestamp 1666464484
transform 1 0 18952 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_206
timestamp 1666464484
transform 1 0 20056 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_218
timestamp 1666464484
transform 1 0 21160 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_230
timestamp 1666464484
transform 1 0 22264 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_237
timestamp 1666464484
transform 1 0 22908 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_249
timestamp 1666464484
transform 1 0 24012 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_261
timestamp 1666464484
transform 1 0 25116 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_273
timestamp 1666464484
transform 1 0 26220 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_280
timestamp 1666464484
transform 1 0 26864 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_292
timestamp 1666464484
transform 1 0 27968 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_304
timestamp 1666464484
transform 1 0 29072 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_316
timestamp 1666464484
transform 1 0 30176 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_323
timestamp 1666464484
transform 1 0 30820 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_335
timestamp 1666464484
transform 1 0 31924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_347
timestamp 1666464484
transform 1 0 33028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_359
timestamp 1666464484
transform 1 0 34132 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_366
timestamp 1666464484
transform 1 0 34776 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_378
timestamp 1666464484
transform 1 0 35880 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_390
timestamp 1666464484
transform 1 0 36984 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_402
timestamp 1666464484
transform 1 0 38088 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_409
timestamp 1666464484
transform 1 0 38732 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1666464484
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1666464484
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_445
timestamp 1666464484
transform 1 0 42044 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_452
timestamp 1666464484
transform 1 0 42688 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_464
timestamp 1666464484
transform 1 0 43792 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_476
timestamp 1666464484
transform 1 0 44896 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_488
timestamp 1666464484
transform 1 0 46000 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_495
timestamp 1666464484
transform 1 0 46644 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_507
timestamp 1666464484
transform 1 0 47748 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_519
timestamp 1666464484
transform 1 0 48852 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_531
timestamp 1666464484
transform 1 0 49956 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_538
timestamp 1666464484
transform 1 0 50600 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_550
timestamp 1666464484
transform 1 0 51704 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_562
timestamp 1666464484
transform 1 0 52808 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_574
timestamp 1666464484
transform 1 0 53912 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_581
timestamp 1666464484
transform 1 0 54556 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_593
timestamp 1666464484
transform 1 0 55660 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_605
timestamp 1666464484
transform 1 0 56764 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_617
timestamp 1666464484
transform 1 0 57868 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_624
timestamp 1666464484
transform 1 0 58512 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666464484
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1666464484
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_39
timestamp 1666464484
transform 1 0 4692 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_44
timestamp 1666464484
transform 1 0 5152 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_56
timestamp 1666464484
transform 1 0 6256 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_68
timestamp 1666464484
transform 1 0 7360 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_80
timestamp 1666464484
transform 1 0 8464 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_87
timestamp 1666464484
transform 1 0 9108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_99
timestamp 1666464484
transform 1 0 10212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_111
timestamp 1666464484
transform 1 0 11316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_123
timestamp 1666464484
transform 1 0 12420 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_130
timestamp 1666464484
transform 1 0 13064 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_142
timestamp 1666464484
transform 1 0 14168 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_154
timestamp 1666464484
transform 1 0 15272 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_166
timestamp 1666464484
transform 1 0 16376 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_173
timestamp 1666464484
transform 1 0 17020 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_185
timestamp 1666464484
transform 1 0 18124 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_197
timestamp 1666464484
transform 1 0 19228 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_209
timestamp 1666464484
transform 1 0 20332 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_216
timestamp 1666464484
transform 1 0 20976 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_228
timestamp 1666464484
transform 1 0 22080 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_240
timestamp 1666464484
transform 1 0 23184 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_252
timestamp 1666464484
transform 1 0 24288 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_259
timestamp 1666464484
transform 1 0 24932 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_271
timestamp 1666464484
transform 1 0 26036 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_283
timestamp 1666464484
transform 1 0 27140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_295
timestamp 1666464484
transform 1 0 28244 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_302
timestamp 1666464484
transform 1 0 28888 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_314
timestamp 1666464484
transform 1 0 29992 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_326
timestamp 1666464484
transform 1 0 31096 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_338
timestamp 1666464484
transform 1 0 32200 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_345
timestamp 1666464484
transform 1 0 32844 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_357
timestamp 1666464484
transform 1 0 33948 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_369
timestamp 1666464484
transform 1 0 35052 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_381
timestamp 1666464484
transform 1 0 36156 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_388
timestamp 1666464484
transform 1 0 36800 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_400
timestamp 1666464484
transform 1 0 37904 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_412
timestamp 1666464484
transform 1 0 39008 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_424
timestamp 1666464484
transform 1 0 40112 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_431
timestamp 1666464484
transform 1 0 40756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_443
timestamp 1666464484
transform 1 0 41860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_455
timestamp 1666464484
transform 1 0 42964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_467
timestamp 1666464484
transform 1 0 44068 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_474
timestamp 1666464484
transform 1 0 44712 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_486
timestamp 1666464484
transform 1 0 45816 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_498
timestamp 1666464484
transform 1 0 46920 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_510
timestamp 1666464484
transform 1 0 48024 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1666464484
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1666464484
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1666464484
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1666464484
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_560
timestamp 1666464484
transform 1 0 52624 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_572
timestamp 1666464484
transform 1 0 53728 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_584
timestamp 1666464484
transform 1 0 54832 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_596
timestamp 1666464484
transform 1 0 55936 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_603
timestamp 1666464484
transform 1 0 56580 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_615
timestamp 1666464484
transform 1 0 57684 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_623
timestamp 1666464484
transform 1 0 58420 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_15
timestamp 1666464484
transform 1 0 2484 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_22
timestamp 1666464484
transform 1 0 3128 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_34
timestamp 1666464484
transform 1 0 4232 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_46
timestamp 1666464484
transform 1 0 5336 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_58
timestamp 1666464484
transform 1 0 6440 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1666464484
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_77
timestamp 1666464484
transform 1 0 8188 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_89
timestamp 1666464484
transform 1 0 9292 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_101
timestamp 1666464484
transform 1 0 10396 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_108
timestamp 1666464484
transform 1 0 11040 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_120
timestamp 1666464484
transform 1 0 12144 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_132
timestamp 1666464484
transform 1 0 13248 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_144
timestamp 1666464484
transform 1 0 14352 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_151
timestamp 1666464484
transform 1 0 14996 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_163
timestamp 1666464484
transform 1 0 16100 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_175
timestamp 1666464484
transform 1 0 17204 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_187
timestamp 1666464484
transform 1 0 18308 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_194
timestamp 1666464484
transform 1 0 18952 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_206
timestamp 1666464484
transform 1 0 20056 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_218
timestamp 1666464484
transform 1 0 21160 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_230
timestamp 1666464484
transform 1 0 22264 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1666464484
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_249
timestamp 1666464484
transform 1 0 24012 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_261
timestamp 1666464484
transform 1 0 25116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_273
timestamp 1666464484
transform 1 0 26220 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_280
timestamp 1666464484
transform 1 0 26864 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_292
timestamp 1666464484
transform 1 0 27968 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_304
timestamp 1666464484
transform 1 0 29072 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_316
timestamp 1666464484
transform 1 0 30176 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_323
timestamp 1666464484
transform 1 0 30820 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_335
timestamp 1666464484
transform 1 0 31924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_347
timestamp 1666464484
transform 1 0 33028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_359
timestamp 1666464484
transform 1 0 34132 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_366
timestamp 1666464484
transform 1 0 34776 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_378
timestamp 1666464484
transform 1 0 35880 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_390
timestamp 1666464484
transform 1 0 36984 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_402
timestamp 1666464484
transform 1 0 38088 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_409
timestamp 1666464484
transform 1 0 38732 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1666464484
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1666464484
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_445
timestamp 1666464484
transform 1 0 42044 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_452
timestamp 1666464484
transform 1 0 42688 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_464
timestamp 1666464484
transform 1 0 43792 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_476
timestamp 1666464484
transform 1 0 44896 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_488
timestamp 1666464484
transform 1 0 46000 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_495
timestamp 1666464484
transform 1 0 46644 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_507
timestamp 1666464484
transform 1 0 47748 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_519
timestamp 1666464484
transform 1 0 48852 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_531
timestamp 1666464484
transform 1 0 49956 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_538
timestamp 1666464484
transform 1 0 50600 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_550
timestamp 1666464484
transform 1 0 51704 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_562
timestamp 1666464484
transform 1 0 52808 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_574
timestamp 1666464484
transform 1 0 53912 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_581
timestamp 1666464484
transform 1 0 54556 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_593
timestamp 1666464484
transform 1 0 55660 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_605
timestamp 1666464484
transform 1 0 56764 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_617
timestamp 1666464484
transform 1 0 57868 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_624
timestamp 1666464484
transform 1 0 58512 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1666464484
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1666464484
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1666464484
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_39
timestamp 1666464484
transform 1 0 4692 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_44
timestamp 1666464484
transform 1 0 5152 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_56
timestamp 1666464484
transform 1 0 6256 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_68
timestamp 1666464484
transform 1 0 7360 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_80
timestamp 1666464484
transform 1 0 8464 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_87
timestamp 1666464484
transform 1 0 9108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_99
timestamp 1666464484
transform 1 0 10212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_111
timestamp 1666464484
transform 1 0 11316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_123
timestamp 1666464484
transform 1 0 12420 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_130
timestamp 1666464484
transform 1 0 13064 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_142
timestamp 1666464484
transform 1 0 14168 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_154
timestamp 1666464484
transform 1 0 15272 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_166
timestamp 1666464484
transform 1 0 16376 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_173
timestamp 1666464484
transform 1 0 17020 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_185
timestamp 1666464484
transform 1 0 18124 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_197
timestamp 1666464484
transform 1 0 19228 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_209
timestamp 1666464484
transform 1 0 20332 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_216
timestamp 1666464484
transform 1 0 20976 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_228
timestamp 1666464484
transform 1 0 22080 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_240
timestamp 1666464484
transform 1 0 23184 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_252
timestamp 1666464484
transform 1 0 24288 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_259
timestamp 1666464484
transform 1 0 24932 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_271
timestamp 1666464484
transform 1 0 26036 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_283
timestamp 1666464484
transform 1 0 27140 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_295
timestamp 1666464484
transform 1 0 28244 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_302
timestamp 1666464484
transform 1 0 28888 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_314
timestamp 1666464484
transform 1 0 29992 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_326
timestamp 1666464484
transform 1 0 31096 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_338
timestamp 1666464484
transform 1 0 32200 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_345
timestamp 1666464484
transform 1 0 32844 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_357
timestamp 1666464484
transform 1 0 33948 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_369
timestamp 1666464484
transform 1 0 35052 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_381
timestamp 1666464484
transform 1 0 36156 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_388
timestamp 1666464484
transform 1 0 36800 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_400
timestamp 1666464484
transform 1 0 37904 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_412
timestamp 1666464484
transform 1 0 39008 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_424
timestamp 1666464484
transform 1 0 40112 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_431
timestamp 1666464484
transform 1 0 40756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_443
timestamp 1666464484
transform 1 0 41860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_455
timestamp 1666464484
transform 1 0 42964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_467
timestamp 1666464484
transform 1 0 44068 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_474
timestamp 1666464484
transform 1 0 44712 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_486
timestamp 1666464484
transform 1 0 45816 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_498
timestamp 1666464484
transform 1 0 46920 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_510
timestamp 1666464484
transform 1 0 48024 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1666464484
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1666464484
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1666464484
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1666464484
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_560
timestamp 1666464484
transform 1 0 52624 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_572
timestamp 1666464484
transform 1 0 53728 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_584
timestamp 1666464484
transform 1 0 54832 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_596
timestamp 1666464484
transform 1 0 55936 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_603
timestamp 1666464484
transform 1 0 56580 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_615
timestamp 1666464484
transform 1 0 57684 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_623
timestamp 1666464484
transform 1 0 58420 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1666464484
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_15
timestamp 1666464484
transform 1 0 2484 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_22
timestamp 1666464484
transform 1 0 3128 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_34
timestamp 1666464484
transform 1 0 4232 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_46
timestamp 1666464484
transform 1 0 5336 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_58
timestamp 1666464484
transform 1 0 6440 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1666464484
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_77
timestamp 1666464484
transform 1 0 8188 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_89
timestamp 1666464484
transform 1 0 9292 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_101
timestamp 1666464484
transform 1 0 10396 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_108
timestamp 1666464484
transform 1 0 11040 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_120
timestamp 1666464484
transform 1 0 12144 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_132
timestamp 1666464484
transform 1 0 13248 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_144
timestamp 1666464484
transform 1 0 14352 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_151
timestamp 1666464484
transform 1 0 14996 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_163
timestamp 1666464484
transform 1 0 16100 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_175
timestamp 1666464484
transform 1 0 17204 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_187
timestamp 1666464484
transform 1 0 18308 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_194
timestamp 1666464484
transform 1 0 18952 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_206
timestamp 1666464484
transform 1 0 20056 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_218
timestamp 1666464484
transform 1 0 21160 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_230
timestamp 1666464484
transform 1 0 22264 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_237
timestamp 1666464484
transform 1 0 22908 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_249
timestamp 1666464484
transform 1 0 24012 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_261
timestamp 1666464484
transform 1 0 25116 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_273
timestamp 1666464484
transform 1 0 26220 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_280
timestamp 1666464484
transform 1 0 26864 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_292
timestamp 1666464484
transform 1 0 27968 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_304
timestamp 1666464484
transform 1 0 29072 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_316
timestamp 1666464484
transform 1 0 30176 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_323
timestamp 1666464484
transform 1 0 30820 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_335
timestamp 1666464484
transform 1 0 31924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_347
timestamp 1666464484
transform 1 0 33028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_359
timestamp 1666464484
transform 1 0 34132 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_366
timestamp 1666464484
transform 1 0 34776 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_378
timestamp 1666464484
transform 1 0 35880 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_390
timestamp 1666464484
transform 1 0 36984 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_402
timestamp 1666464484
transform 1 0 38088 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_409
timestamp 1666464484
transform 1 0 38732 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1666464484
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1666464484
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_445
timestamp 1666464484
transform 1 0 42044 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_452
timestamp 1666464484
transform 1 0 42688 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_464
timestamp 1666464484
transform 1 0 43792 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_476
timestamp 1666464484
transform 1 0 44896 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_488
timestamp 1666464484
transform 1 0 46000 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_495
timestamp 1666464484
transform 1 0 46644 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_507
timestamp 1666464484
transform 1 0 47748 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_519
timestamp 1666464484
transform 1 0 48852 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_531
timestamp 1666464484
transform 1 0 49956 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_538
timestamp 1666464484
transform 1 0 50600 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_550
timestamp 1666464484
transform 1 0 51704 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_562
timestamp 1666464484
transform 1 0 52808 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_574
timestamp 1666464484
transform 1 0 53912 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_581
timestamp 1666464484
transform 1 0 54556 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_593
timestamp 1666464484
transform 1 0 55660 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_605
timestamp 1666464484
transform 1 0 56764 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_617
timestamp 1666464484
transform 1 0 57868 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_624
timestamp 1666464484
transform 1 0 58512 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1666464484
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1666464484
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1666464484
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_39
timestamp 1666464484
transform 1 0 4692 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_44
timestamp 1666464484
transform 1 0 5152 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_56
timestamp 1666464484
transform 1 0 6256 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_68
timestamp 1666464484
transform 1 0 7360 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_80
timestamp 1666464484
transform 1 0 8464 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_87
timestamp 1666464484
transform 1 0 9108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_99
timestamp 1666464484
transform 1 0 10212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_111
timestamp 1666464484
transform 1 0 11316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_123
timestamp 1666464484
transform 1 0 12420 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_130
timestamp 1666464484
transform 1 0 13064 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_142
timestamp 1666464484
transform 1 0 14168 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_154
timestamp 1666464484
transform 1 0 15272 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_166
timestamp 1666464484
transform 1 0 16376 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_173
timestamp 1666464484
transform 1 0 17020 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_185
timestamp 1666464484
transform 1 0 18124 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_197
timestamp 1666464484
transform 1 0 19228 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_209
timestamp 1666464484
transform 1 0 20332 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_216
timestamp 1666464484
transform 1 0 20976 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_228
timestamp 1666464484
transform 1 0 22080 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_240
timestamp 1666464484
transform 1 0 23184 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_252
timestamp 1666464484
transform 1 0 24288 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_259
timestamp 1666464484
transform 1 0 24932 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_271
timestamp 1666464484
transform 1 0 26036 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_283
timestamp 1666464484
transform 1 0 27140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_295
timestamp 1666464484
transform 1 0 28244 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_302
timestamp 1666464484
transform 1 0 28888 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_314
timestamp 1666464484
transform 1 0 29992 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_326
timestamp 1666464484
transform 1 0 31096 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_338
timestamp 1666464484
transform 1 0 32200 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_345
timestamp 1666464484
transform 1 0 32844 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_357
timestamp 1666464484
transform 1 0 33948 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_369
timestamp 1666464484
transform 1 0 35052 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_381
timestamp 1666464484
transform 1 0 36156 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_388
timestamp 1666464484
transform 1 0 36800 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_400
timestamp 1666464484
transform 1 0 37904 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_412
timestamp 1666464484
transform 1 0 39008 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_424
timestamp 1666464484
transform 1 0 40112 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_431
timestamp 1666464484
transform 1 0 40756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_443
timestamp 1666464484
transform 1 0 41860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_455
timestamp 1666464484
transform 1 0 42964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_467
timestamp 1666464484
transform 1 0 44068 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_474
timestamp 1666464484
transform 1 0 44712 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_486
timestamp 1666464484
transform 1 0 45816 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_498
timestamp 1666464484
transform 1 0 46920 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_510
timestamp 1666464484
transform 1 0 48024 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1666464484
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1666464484
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1666464484
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1666464484
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_560
timestamp 1666464484
transform 1 0 52624 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_572
timestamp 1666464484
transform 1 0 53728 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_584
timestamp 1666464484
transform 1 0 54832 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_596
timestamp 1666464484
transform 1 0 55936 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_603
timestamp 1666464484
transform 1 0 56580 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_615
timestamp 1666464484
transform 1 0 57684 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_623
timestamp 1666464484
transform 1 0 58420 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1666464484
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_15
timestamp 1666464484
transform 1 0 2484 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_22
timestamp 1666464484
transform 1 0 3128 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_34
timestamp 1666464484
transform 1 0 4232 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_46
timestamp 1666464484
transform 1 0 5336 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_58
timestamp 1666464484
transform 1 0 6440 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1666464484
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_77
timestamp 1666464484
transform 1 0 8188 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_89
timestamp 1666464484
transform 1 0 9292 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_101
timestamp 1666464484
transform 1 0 10396 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_108
timestamp 1666464484
transform 1 0 11040 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_120
timestamp 1666464484
transform 1 0 12144 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_132
timestamp 1666464484
transform 1 0 13248 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_144
timestamp 1666464484
transform 1 0 14352 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_151
timestamp 1666464484
transform 1 0 14996 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_163
timestamp 1666464484
transform 1 0 16100 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_175
timestamp 1666464484
transform 1 0 17204 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_187
timestamp 1666464484
transform 1 0 18308 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_194
timestamp 1666464484
transform 1 0 18952 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_206
timestamp 1666464484
transform 1 0 20056 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_218
timestamp 1666464484
transform 1 0 21160 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_230
timestamp 1666464484
transform 1 0 22264 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_237
timestamp 1666464484
transform 1 0 22908 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_249
timestamp 1666464484
transform 1 0 24012 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_261
timestamp 1666464484
transform 1 0 25116 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_273
timestamp 1666464484
transform 1 0 26220 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_280
timestamp 1666464484
transform 1 0 26864 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_292
timestamp 1666464484
transform 1 0 27968 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_304
timestamp 1666464484
transform 1 0 29072 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_316
timestamp 1666464484
transform 1 0 30176 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_323
timestamp 1666464484
transform 1 0 30820 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_335
timestamp 1666464484
transform 1 0 31924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_347
timestamp 1666464484
transform 1 0 33028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_359
timestamp 1666464484
transform 1 0 34132 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_366
timestamp 1666464484
transform 1 0 34776 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_378
timestamp 1666464484
transform 1 0 35880 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_390
timestamp 1666464484
transform 1 0 36984 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_402
timestamp 1666464484
transform 1 0 38088 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_409
timestamp 1666464484
transform 1 0 38732 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1666464484
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1666464484
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_445
timestamp 1666464484
transform 1 0 42044 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_452
timestamp 1666464484
transform 1 0 42688 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_464
timestamp 1666464484
transform 1 0 43792 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_476
timestamp 1666464484
transform 1 0 44896 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_488
timestamp 1666464484
transform 1 0 46000 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_495
timestamp 1666464484
transform 1 0 46644 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_507
timestamp 1666464484
transform 1 0 47748 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_519
timestamp 1666464484
transform 1 0 48852 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_531
timestamp 1666464484
transform 1 0 49956 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_538
timestamp 1666464484
transform 1 0 50600 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_550
timestamp 1666464484
transform 1 0 51704 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_562
timestamp 1666464484
transform 1 0 52808 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_574
timestamp 1666464484
transform 1 0 53912 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_581
timestamp 1666464484
transform 1 0 54556 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_593
timestamp 1666464484
transform 1 0 55660 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_605
timestamp 1666464484
transform 1 0 56764 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_617
timestamp 1666464484
transform 1 0 57868 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_624
timestamp 1666464484
transform 1 0 58512 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1666464484
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1666464484
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1666464484
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_39
timestamp 1666464484
transform 1 0 4692 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_44
timestamp 1666464484
transform 1 0 5152 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_56
timestamp 1666464484
transform 1 0 6256 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_68
timestamp 1666464484
transform 1 0 7360 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_80
timestamp 1666464484
transform 1 0 8464 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_87
timestamp 1666464484
transform 1 0 9108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_99
timestamp 1666464484
transform 1 0 10212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_111
timestamp 1666464484
transform 1 0 11316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_123
timestamp 1666464484
transform 1 0 12420 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_130
timestamp 1666464484
transform 1 0 13064 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_142
timestamp 1666464484
transform 1 0 14168 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_154
timestamp 1666464484
transform 1 0 15272 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_166
timestamp 1666464484
transform 1 0 16376 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_173
timestamp 1666464484
transform 1 0 17020 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_185
timestamp 1666464484
transform 1 0 18124 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_197
timestamp 1666464484
transform 1 0 19228 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_209
timestamp 1666464484
transform 1 0 20332 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_216
timestamp 1666464484
transform 1 0 20976 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_228
timestamp 1666464484
transform 1 0 22080 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_240
timestamp 1666464484
transform 1 0 23184 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_252
timestamp 1666464484
transform 1 0 24288 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_259
timestamp 1666464484
transform 1 0 24932 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_271
timestamp 1666464484
transform 1 0 26036 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_283
timestamp 1666464484
transform 1 0 27140 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_295
timestamp 1666464484
transform 1 0 28244 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_302
timestamp 1666464484
transform 1 0 28888 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_314
timestamp 1666464484
transform 1 0 29992 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_326
timestamp 1666464484
transform 1 0 31096 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_338
timestamp 1666464484
transform 1 0 32200 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_345
timestamp 1666464484
transform 1 0 32844 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_357
timestamp 1666464484
transform 1 0 33948 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_369
timestamp 1666464484
transform 1 0 35052 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_381
timestamp 1666464484
transform 1 0 36156 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_388
timestamp 1666464484
transform 1 0 36800 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_400
timestamp 1666464484
transform 1 0 37904 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_412
timestamp 1666464484
transform 1 0 39008 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_424
timestamp 1666464484
transform 1 0 40112 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_431
timestamp 1666464484
transform 1 0 40756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_443
timestamp 1666464484
transform 1 0 41860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_455
timestamp 1666464484
transform 1 0 42964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_467
timestamp 1666464484
transform 1 0 44068 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_474
timestamp 1666464484
transform 1 0 44712 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_486
timestamp 1666464484
transform 1 0 45816 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_498
timestamp 1666464484
transform 1 0 46920 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_510
timestamp 1666464484
transform 1 0 48024 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1666464484
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1666464484
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1666464484
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1666464484
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_560
timestamp 1666464484
transform 1 0 52624 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_572
timestamp 1666464484
transform 1 0 53728 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_584
timestamp 1666464484
transform 1 0 54832 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_596
timestamp 1666464484
transform 1 0 55936 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_603
timestamp 1666464484
transform 1 0 56580 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_615
timestamp 1666464484
transform 1 0 57684 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_623
timestamp 1666464484
transform 1 0 58420 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1666464484
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_15
timestamp 1666464484
transform 1 0 2484 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_22
timestamp 1666464484
transform 1 0 3128 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_34
timestamp 1666464484
transform 1 0 4232 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_46
timestamp 1666464484
transform 1 0 5336 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_58
timestamp 1666464484
transform 1 0 6440 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1666464484
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_77
timestamp 1666464484
transform 1 0 8188 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_89
timestamp 1666464484
transform 1 0 9292 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_101
timestamp 1666464484
transform 1 0 10396 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_108
timestamp 1666464484
transform 1 0 11040 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_120
timestamp 1666464484
transform 1 0 12144 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_132
timestamp 1666464484
transform 1 0 13248 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_144
timestamp 1666464484
transform 1 0 14352 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_151
timestamp 1666464484
transform 1 0 14996 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_163
timestamp 1666464484
transform 1 0 16100 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_175
timestamp 1666464484
transform 1 0 17204 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_187
timestamp 1666464484
transform 1 0 18308 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_194
timestamp 1666464484
transform 1 0 18952 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_206
timestamp 1666464484
transform 1 0 20056 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_218
timestamp 1666464484
transform 1 0 21160 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_230
timestamp 1666464484
transform 1 0 22264 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_237
timestamp 1666464484
transform 1 0 22908 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_249
timestamp 1666464484
transform 1 0 24012 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_261
timestamp 1666464484
transform 1 0 25116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_273
timestamp 1666464484
transform 1 0 26220 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_280
timestamp 1666464484
transform 1 0 26864 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_292
timestamp 1666464484
transform 1 0 27968 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_304
timestamp 1666464484
transform 1 0 29072 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_316
timestamp 1666464484
transform 1 0 30176 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_323
timestamp 1666464484
transform 1 0 30820 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_335
timestamp 1666464484
transform 1 0 31924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_347
timestamp 1666464484
transform 1 0 33028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_359
timestamp 1666464484
transform 1 0 34132 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_366
timestamp 1666464484
transform 1 0 34776 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_378
timestamp 1666464484
transform 1 0 35880 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_390
timestamp 1666464484
transform 1 0 36984 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_402
timestamp 1666464484
transform 1 0 38088 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_409
timestamp 1666464484
transform 1 0 38732 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1666464484
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1666464484
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_445
timestamp 1666464484
transform 1 0 42044 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_452
timestamp 1666464484
transform 1 0 42688 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_464
timestamp 1666464484
transform 1 0 43792 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_476
timestamp 1666464484
transform 1 0 44896 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_488
timestamp 1666464484
transform 1 0 46000 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_495
timestamp 1666464484
transform 1 0 46644 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_507
timestamp 1666464484
transform 1 0 47748 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_519
timestamp 1666464484
transform 1 0 48852 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_531
timestamp 1666464484
transform 1 0 49956 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_538
timestamp 1666464484
transform 1 0 50600 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_550
timestamp 1666464484
transform 1 0 51704 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_562
timestamp 1666464484
transform 1 0 52808 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_574
timestamp 1666464484
transform 1 0 53912 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_581
timestamp 1666464484
transform 1 0 54556 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_593
timestamp 1666464484
transform 1 0 55660 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_605
timestamp 1666464484
transform 1 0 56764 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_617
timestamp 1666464484
transform 1 0 57868 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_624
timestamp 1666464484
transform 1 0 58512 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1666464484
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1666464484
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1666464484
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_39
timestamp 1666464484
transform 1 0 4692 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_44
timestamp 1666464484
transform 1 0 5152 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_56
timestamp 1666464484
transform 1 0 6256 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_68
timestamp 1666464484
transform 1 0 7360 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_80
timestamp 1666464484
transform 1 0 8464 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_87
timestamp 1666464484
transform 1 0 9108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_99
timestamp 1666464484
transform 1 0 10212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_111
timestamp 1666464484
transform 1 0 11316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_123
timestamp 1666464484
transform 1 0 12420 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_130
timestamp 1666464484
transform 1 0 13064 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_142
timestamp 1666464484
transform 1 0 14168 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_154
timestamp 1666464484
transform 1 0 15272 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_166
timestamp 1666464484
transform 1 0 16376 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_173
timestamp 1666464484
transform 1 0 17020 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_185
timestamp 1666464484
transform 1 0 18124 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_197
timestamp 1666464484
transform 1 0 19228 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_209
timestamp 1666464484
transform 1 0 20332 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_216
timestamp 1666464484
transform 1 0 20976 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_228
timestamp 1666464484
transform 1 0 22080 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_240
timestamp 1666464484
transform 1 0 23184 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_252
timestamp 1666464484
transform 1 0 24288 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_259
timestamp 1666464484
transform 1 0 24932 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_271
timestamp 1666464484
transform 1 0 26036 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_283
timestamp 1666464484
transform 1 0 27140 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_295
timestamp 1666464484
transform 1 0 28244 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_302
timestamp 1666464484
transform 1 0 28888 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_314
timestamp 1666464484
transform 1 0 29992 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_326
timestamp 1666464484
transform 1 0 31096 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_338
timestamp 1666464484
transform 1 0 32200 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_345
timestamp 1666464484
transform 1 0 32844 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_357
timestamp 1666464484
transform 1 0 33948 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_369
timestamp 1666464484
transform 1 0 35052 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_381
timestamp 1666464484
transform 1 0 36156 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_388
timestamp 1666464484
transform 1 0 36800 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_400
timestamp 1666464484
transform 1 0 37904 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_412
timestamp 1666464484
transform 1 0 39008 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_424
timestamp 1666464484
transform 1 0 40112 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_431
timestamp 1666464484
transform 1 0 40756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_443
timestamp 1666464484
transform 1 0 41860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_455
timestamp 1666464484
transform 1 0 42964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_467
timestamp 1666464484
transform 1 0 44068 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_474
timestamp 1666464484
transform 1 0 44712 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_486
timestamp 1666464484
transform 1 0 45816 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_498
timestamp 1666464484
transform 1 0 46920 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_510
timestamp 1666464484
transform 1 0 48024 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1666464484
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1666464484
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1666464484
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1666464484
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_560
timestamp 1666464484
transform 1 0 52624 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_572
timestamp 1666464484
transform 1 0 53728 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_584
timestamp 1666464484
transform 1 0 54832 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_596
timestamp 1666464484
transform 1 0 55936 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_603
timestamp 1666464484
transform 1 0 56580 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_615
timestamp 1666464484
transform 1 0 57684 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_623
timestamp 1666464484
transform 1 0 58420 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1666464484
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_15
timestamp 1666464484
transform 1 0 2484 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_22
timestamp 1666464484
transform 1 0 3128 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_34
timestamp 1666464484
transform 1 0 4232 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_46
timestamp 1666464484
transform 1 0 5336 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_58
timestamp 1666464484
transform 1 0 6440 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1666464484
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_77
timestamp 1666464484
transform 1 0 8188 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_89
timestamp 1666464484
transform 1 0 9292 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_101
timestamp 1666464484
transform 1 0 10396 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_108
timestamp 1666464484
transform 1 0 11040 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_120
timestamp 1666464484
transform 1 0 12144 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_132
timestamp 1666464484
transform 1 0 13248 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_144
timestamp 1666464484
transform 1 0 14352 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_151
timestamp 1666464484
transform 1 0 14996 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_163
timestamp 1666464484
transform 1 0 16100 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_175
timestamp 1666464484
transform 1 0 17204 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_187
timestamp 1666464484
transform 1 0 18308 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_194
timestamp 1666464484
transform 1 0 18952 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_206
timestamp 1666464484
transform 1 0 20056 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_218
timestamp 1666464484
transform 1 0 21160 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_230
timestamp 1666464484
transform 1 0 22264 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_237
timestamp 1666464484
transform 1 0 22908 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_249
timestamp 1666464484
transform 1 0 24012 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_261
timestamp 1666464484
transform 1 0 25116 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_273
timestamp 1666464484
transform 1 0 26220 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_280
timestamp 1666464484
transform 1 0 26864 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_292
timestamp 1666464484
transform 1 0 27968 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_304
timestamp 1666464484
transform 1 0 29072 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_316
timestamp 1666464484
transform 1 0 30176 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_323
timestamp 1666464484
transform 1 0 30820 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_335
timestamp 1666464484
transform 1 0 31924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_347
timestamp 1666464484
transform 1 0 33028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_359
timestamp 1666464484
transform 1 0 34132 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_366
timestamp 1666464484
transform 1 0 34776 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_378
timestamp 1666464484
transform 1 0 35880 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_390
timestamp 1666464484
transform 1 0 36984 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_402
timestamp 1666464484
transform 1 0 38088 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_409
timestamp 1666464484
transform 1 0 38732 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1666464484
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1666464484
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_445
timestamp 1666464484
transform 1 0 42044 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_452
timestamp 1666464484
transform 1 0 42688 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_464
timestamp 1666464484
transform 1 0 43792 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_476
timestamp 1666464484
transform 1 0 44896 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_488
timestamp 1666464484
transform 1 0 46000 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_495
timestamp 1666464484
transform 1 0 46644 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_507
timestamp 1666464484
transform 1 0 47748 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_519
timestamp 1666464484
transform 1 0 48852 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_531
timestamp 1666464484
transform 1 0 49956 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_538
timestamp 1666464484
transform 1 0 50600 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_550
timestamp 1666464484
transform 1 0 51704 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_562
timestamp 1666464484
transform 1 0 52808 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_574
timestamp 1666464484
transform 1 0 53912 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_581
timestamp 1666464484
transform 1 0 54556 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_593
timestamp 1666464484
transform 1 0 55660 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_605
timestamp 1666464484
transform 1 0 56764 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_617
timestamp 1666464484
transform 1 0 57868 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_624
timestamp 1666464484
transform 1 0 58512 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1666464484
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1666464484
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1666464484
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_39
timestamp 1666464484
transform 1 0 4692 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_44
timestamp 1666464484
transform 1 0 5152 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_56
timestamp 1666464484
transform 1 0 6256 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_68
timestamp 1666464484
transform 1 0 7360 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_80
timestamp 1666464484
transform 1 0 8464 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_87
timestamp 1666464484
transform 1 0 9108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_99
timestamp 1666464484
transform 1 0 10212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_111
timestamp 1666464484
transform 1 0 11316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_123
timestamp 1666464484
transform 1 0 12420 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_130
timestamp 1666464484
transform 1 0 13064 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_142
timestamp 1666464484
transform 1 0 14168 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_154
timestamp 1666464484
transform 1 0 15272 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_166
timestamp 1666464484
transform 1 0 16376 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_173
timestamp 1666464484
transform 1 0 17020 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_185
timestamp 1666464484
transform 1 0 18124 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_197
timestamp 1666464484
transform 1 0 19228 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_209
timestamp 1666464484
transform 1 0 20332 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_216
timestamp 1666464484
transform 1 0 20976 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_228
timestamp 1666464484
transform 1 0 22080 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_240
timestamp 1666464484
transform 1 0 23184 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_252
timestamp 1666464484
transform 1 0 24288 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_259
timestamp 1666464484
transform 1 0 24932 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_271
timestamp 1666464484
transform 1 0 26036 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_283
timestamp 1666464484
transform 1 0 27140 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_295
timestamp 1666464484
transform 1 0 28244 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_302
timestamp 1666464484
transform 1 0 28888 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_314
timestamp 1666464484
transform 1 0 29992 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_326
timestamp 1666464484
transform 1 0 31096 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_338
timestamp 1666464484
transform 1 0 32200 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_345
timestamp 1666464484
transform 1 0 32844 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_357
timestamp 1666464484
transform 1 0 33948 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_369
timestamp 1666464484
transform 1 0 35052 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_381
timestamp 1666464484
transform 1 0 36156 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_388
timestamp 1666464484
transform 1 0 36800 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_400
timestamp 1666464484
transform 1 0 37904 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_412
timestamp 1666464484
transform 1 0 39008 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_424
timestamp 1666464484
transform 1 0 40112 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_431
timestamp 1666464484
transform 1 0 40756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_443
timestamp 1666464484
transform 1 0 41860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_455
timestamp 1666464484
transform 1 0 42964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_467
timestamp 1666464484
transform 1 0 44068 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_474
timestamp 1666464484
transform 1 0 44712 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_486
timestamp 1666464484
transform 1 0 45816 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_498
timestamp 1666464484
transform 1 0 46920 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_510
timestamp 1666464484
transform 1 0 48024 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1666464484
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1666464484
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1666464484
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1666464484
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_560
timestamp 1666464484
transform 1 0 52624 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_572
timestamp 1666464484
transform 1 0 53728 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_584
timestamp 1666464484
transform 1 0 54832 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_596
timestamp 1666464484
transform 1 0 55936 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_603
timestamp 1666464484
transform 1 0 56580 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_615
timestamp 1666464484
transform 1 0 57684 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_623
timestamp 1666464484
transform 1 0 58420 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1666464484
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_15
timestamp 1666464484
transform 1 0 2484 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_22
timestamp 1666464484
transform 1 0 3128 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_34
timestamp 1666464484
transform 1 0 4232 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_46
timestamp 1666464484
transform 1 0 5336 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_58
timestamp 1666464484
transform 1 0 6440 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1666464484
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_77
timestamp 1666464484
transform 1 0 8188 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_89
timestamp 1666464484
transform 1 0 9292 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_101
timestamp 1666464484
transform 1 0 10396 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_108
timestamp 1666464484
transform 1 0 11040 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_120
timestamp 1666464484
transform 1 0 12144 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_132
timestamp 1666464484
transform 1 0 13248 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_144
timestamp 1666464484
transform 1 0 14352 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_151
timestamp 1666464484
transform 1 0 14996 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_163
timestamp 1666464484
transform 1 0 16100 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_175
timestamp 1666464484
transform 1 0 17204 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_187
timestamp 1666464484
transform 1 0 18308 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_194
timestamp 1666464484
transform 1 0 18952 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_206
timestamp 1666464484
transform 1 0 20056 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_218
timestamp 1666464484
transform 1 0 21160 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_230
timestamp 1666464484
transform 1 0 22264 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_237
timestamp 1666464484
transform 1 0 22908 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_249
timestamp 1666464484
transform 1 0 24012 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_261
timestamp 1666464484
transform 1 0 25116 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_273
timestamp 1666464484
transform 1 0 26220 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_280
timestamp 1666464484
transform 1 0 26864 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_292
timestamp 1666464484
transform 1 0 27968 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_304
timestamp 1666464484
transform 1 0 29072 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_316
timestamp 1666464484
transform 1 0 30176 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_323
timestamp 1666464484
transform 1 0 30820 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_335
timestamp 1666464484
transform 1 0 31924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_347
timestamp 1666464484
transform 1 0 33028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_359
timestamp 1666464484
transform 1 0 34132 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_366
timestamp 1666464484
transform 1 0 34776 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_378
timestamp 1666464484
transform 1 0 35880 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_390
timestamp 1666464484
transform 1 0 36984 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_402
timestamp 1666464484
transform 1 0 38088 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_409
timestamp 1666464484
transform 1 0 38732 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1666464484
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1666464484
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_445
timestamp 1666464484
transform 1 0 42044 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_452
timestamp 1666464484
transform 1 0 42688 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_464
timestamp 1666464484
transform 1 0 43792 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_476
timestamp 1666464484
transform 1 0 44896 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_488
timestamp 1666464484
transform 1 0 46000 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_495
timestamp 1666464484
transform 1 0 46644 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_507
timestamp 1666464484
transform 1 0 47748 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_519
timestamp 1666464484
transform 1 0 48852 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_531
timestamp 1666464484
transform 1 0 49956 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_538
timestamp 1666464484
transform 1 0 50600 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_550
timestamp 1666464484
transform 1 0 51704 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_562
timestamp 1666464484
transform 1 0 52808 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_574
timestamp 1666464484
transform 1 0 53912 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_581
timestamp 1666464484
transform 1 0 54556 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_593
timestamp 1666464484
transform 1 0 55660 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_605
timestamp 1666464484
transform 1 0 56764 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_617
timestamp 1666464484
transform 1 0 57868 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_624
timestamp 1666464484
transform 1 0 58512 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1666464484
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1666464484
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1666464484
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_39
timestamp 1666464484
transform 1 0 4692 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_44
timestamp 1666464484
transform 1 0 5152 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_56
timestamp 1666464484
transform 1 0 6256 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_68
timestamp 1666464484
transform 1 0 7360 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_80
timestamp 1666464484
transform 1 0 8464 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_87
timestamp 1666464484
transform 1 0 9108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_99
timestamp 1666464484
transform 1 0 10212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_111
timestamp 1666464484
transform 1 0 11316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_123
timestamp 1666464484
transform 1 0 12420 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_130
timestamp 1666464484
transform 1 0 13064 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_142
timestamp 1666464484
transform 1 0 14168 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_154
timestamp 1666464484
transform 1 0 15272 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_166
timestamp 1666464484
transform 1 0 16376 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_173
timestamp 1666464484
transform 1 0 17020 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_185
timestamp 1666464484
transform 1 0 18124 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_197
timestamp 1666464484
transform 1 0 19228 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_209
timestamp 1666464484
transform 1 0 20332 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_216
timestamp 1666464484
transform 1 0 20976 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_228
timestamp 1666464484
transform 1 0 22080 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_240
timestamp 1666464484
transform 1 0 23184 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_252
timestamp 1666464484
transform 1 0 24288 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_259
timestamp 1666464484
transform 1 0 24932 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_271
timestamp 1666464484
transform 1 0 26036 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_283
timestamp 1666464484
transform 1 0 27140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_295
timestamp 1666464484
transform 1 0 28244 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_302
timestamp 1666464484
transform 1 0 28888 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_314
timestamp 1666464484
transform 1 0 29992 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_326
timestamp 1666464484
transform 1 0 31096 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_338
timestamp 1666464484
transform 1 0 32200 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_345
timestamp 1666464484
transform 1 0 32844 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_357
timestamp 1666464484
transform 1 0 33948 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_369
timestamp 1666464484
transform 1 0 35052 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_381
timestamp 1666464484
transform 1 0 36156 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_388
timestamp 1666464484
transform 1 0 36800 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_400
timestamp 1666464484
transform 1 0 37904 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_412
timestamp 1666464484
transform 1 0 39008 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_424
timestamp 1666464484
transform 1 0 40112 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_431
timestamp 1666464484
transform 1 0 40756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_443
timestamp 1666464484
transform 1 0 41860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_455
timestamp 1666464484
transform 1 0 42964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_467
timestamp 1666464484
transform 1 0 44068 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_474
timestamp 1666464484
transform 1 0 44712 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_486
timestamp 1666464484
transform 1 0 45816 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_498
timestamp 1666464484
transform 1 0 46920 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_510
timestamp 1666464484
transform 1 0 48024 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1666464484
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1666464484
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1666464484
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1666464484
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_560
timestamp 1666464484
transform 1 0 52624 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_572
timestamp 1666464484
transform 1 0 53728 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_584
timestamp 1666464484
transform 1 0 54832 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_596
timestamp 1666464484
transform 1 0 55936 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_603
timestamp 1666464484
transform 1 0 56580 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_615
timestamp 1666464484
transform 1 0 57684 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_623
timestamp 1666464484
transform 1 0 58420 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1666464484
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_15
timestamp 1666464484
transform 1 0 2484 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_22
timestamp 1666464484
transform 1 0 3128 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_34
timestamp 1666464484
transform 1 0 4232 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_46
timestamp 1666464484
transform 1 0 5336 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_58
timestamp 1666464484
transform 1 0 6440 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1666464484
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_77
timestamp 1666464484
transform 1 0 8188 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_89
timestamp 1666464484
transform 1 0 9292 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_101
timestamp 1666464484
transform 1 0 10396 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_108
timestamp 1666464484
transform 1 0 11040 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_120
timestamp 1666464484
transform 1 0 12144 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_132
timestamp 1666464484
transform 1 0 13248 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_144
timestamp 1666464484
transform 1 0 14352 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_151
timestamp 1666464484
transform 1 0 14996 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_163
timestamp 1666464484
transform 1 0 16100 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_175
timestamp 1666464484
transform 1 0 17204 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_187
timestamp 1666464484
transform 1 0 18308 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_194
timestamp 1666464484
transform 1 0 18952 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_206
timestamp 1666464484
transform 1 0 20056 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_218
timestamp 1666464484
transform 1 0 21160 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_230
timestamp 1666464484
transform 1 0 22264 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_237
timestamp 1666464484
transform 1 0 22908 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_249
timestamp 1666464484
transform 1 0 24012 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_261
timestamp 1666464484
transform 1 0 25116 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_273
timestamp 1666464484
transform 1 0 26220 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_280
timestamp 1666464484
transform 1 0 26864 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_292
timestamp 1666464484
transform 1 0 27968 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_304
timestamp 1666464484
transform 1 0 29072 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_316
timestamp 1666464484
transform 1 0 30176 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_323
timestamp 1666464484
transform 1 0 30820 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_335
timestamp 1666464484
transform 1 0 31924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_347
timestamp 1666464484
transform 1 0 33028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_359
timestamp 1666464484
transform 1 0 34132 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_366
timestamp 1666464484
transform 1 0 34776 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_378
timestamp 1666464484
transform 1 0 35880 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_390
timestamp 1666464484
transform 1 0 36984 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_402
timestamp 1666464484
transform 1 0 38088 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_409
timestamp 1666464484
transform 1 0 38732 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1666464484
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1666464484
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_445
timestamp 1666464484
transform 1 0 42044 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_452
timestamp 1666464484
transform 1 0 42688 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_464
timestamp 1666464484
transform 1 0 43792 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_476
timestamp 1666464484
transform 1 0 44896 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_488
timestamp 1666464484
transform 1 0 46000 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_495
timestamp 1666464484
transform 1 0 46644 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_507
timestamp 1666464484
transform 1 0 47748 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_519
timestamp 1666464484
transform 1 0 48852 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_531
timestamp 1666464484
transform 1 0 49956 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_538
timestamp 1666464484
transform 1 0 50600 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_550
timestamp 1666464484
transform 1 0 51704 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_562
timestamp 1666464484
transform 1 0 52808 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_574
timestamp 1666464484
transform 1 0 53912 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_581
timestamp 1666464484
transform 1 0 54556 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_593
timestamp 1666464484
transform 1 0 55660 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_605
timestamp 1666464484
transform 1 0 56764 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_617
timestamp 1666464484
transform 1 0 57868 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_624
timestamp 1666464484
transform 1 0 58512 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1666464484
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1666464484
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1666464484
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_39
timestamp 1666464484
transform 1 0 4692 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_44
timestamp 1666464484
transform 1 0 5152 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_56
timestamp 1666464484
transform 1 0 6256 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_68
timestamp 1666464484
transform 1 0 7360 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_80
timestamp 1666464484
transform 1 0 8464 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_87
timestamp 1666464484
transform 1 0 9108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_99
timestamp 1666464484
transform 1 0 10212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_111
timestamp 1666464484
transform 1 0 11316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_123
timestamp 1666464484
transform 1 0 12420 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_130
timestamp 1666464484
transform 1 0 13064 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_142
timestamp 1666464484
transform 1 0 14168 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_154
timestamp 1666464484
transform 1 0 15272 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_166
timestamp 1666464484
transform 1 0 16376 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_173
timestamp 1666464484
transform 1 0 17020 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_185
timestamp 1666464484
transform 1 0 18124 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_197
timestamp 1666464484
transform 1 0 19228 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_209
timestamp 1666464484
transform 1 0 20332 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_216
timestamp 1666464484
transform 1 0 20976 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_228
timestamp 1666464484
transform 1 0 22080 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_240
timestamp 1666464484
transform 1 0 23184 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_252
timestamp 1666464484
transform 1 0 24288 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_259
timestamp 1666464484
transform 1 0 24932 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_271
timestamp 1666464484
transform 1 0 26036 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_283
timestamp 1666464484
transform 1 0 27140 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_295
timestamp 1666464484
transform 1 0 28244 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_302
timestamp 1666464484
transform 1 0 28888 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_314
timestamp 1666464484
transform 1 0 29992 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_326
timestamp 1666464484
transform 1 0 31096 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_338
timestamp 1666464484
transform 1 0 32200 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_345
timestamp 1666464484
transform 1 0 32844 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_357
timestamp 1666464484
transform 1 0 33948 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_369
timestamp 1666464484
transform 1 0 35052 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_381
timestamp 1666464484
transform 1 0 36156 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_388
timestamp 1666464484
transform 1 0 36800 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_400
timestamp 1666464484
transform 1 0 37904 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_412
timestamp 1666464484
transform 1 0 39008 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_424
timestamp 1666464484
transform 1 0 40112 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_431
timestamp 1666464484
transform 1 0 40756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_443
timestamp 1666464484
transform 1 0 41860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_455
timestamp 1666464484
transform 1 0 42964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_467
timestamp 1666464484
transform 1 0 44068 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_474
timestamp 1666464484
transform 1 0 44712 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_486
timestamp 1666464484
transform 1 0 45816 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_498
timestamp 1666464484
transform 1 0 46920 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_510
timestamp 1666464484
transform 1 0 48024 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1666464484
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1666464484
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1666464484
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1666464484
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_560
timestamp 1666464484
transform 1 0 52624 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_572
timestamp 1666464484
transform 1 0 53728 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_584
timestamp 1666464484
transform 1 0 54832 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_596
timestamp 1666464484
transform 1 0 55936 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_603
timestamp 1666464484
transform 1 0 56580 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_615
timestamp 1666464484
transform 1 0 57684 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_623
timestamp 1666464484
transform 1 0 58420 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1666464484
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_15
timestamp 1666464484
transform 1 0 2484 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_22
timestamp 1666464484
transform 1 0 3128 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_34
timestamp 1666464484
transform 1 0 4232 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_46
timestamp 1666464484
transform 1 0 5336 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_58
timestamp 1666464484
transform 1 0 6440 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1666464484
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_77
timestamp 1666464484
transform 1 0 8188 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_89
timestamp 1666464484
transform 1 0 9292 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_101
timestamp 1666464484
transform 1 0 10396 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_108
timestamp 1666464484
transform 1 0 11040 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_120
timestamp 1666464484
transform 1 0 12144 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_132
timestamp 1666464484
transform 1 0 13248 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_144
timestamp 1666464484
transform 1 0 14352 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_151
timestamp 1666464484
transform 1 0 14996 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_163
timestamp 1666464484
transform 1 0 16100 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_175
timestamp 1666464484
transform 1 0 17204 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_187
timestamp 1666464484
transform 1 0 18308 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_194
timestamp 1666464484
transform 1 0 18952 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_206
timestamp 1666464484
transform 1 0 20056 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_218
timestamp 1666464484
transform 1 0 21160 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_230
timestamp 1666464484
transform 1 0 22264 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_237
timestamp 1666464484
transform 1 0 22908 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_249
timestamp 1666464484
transform 1 0 24012 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_261
timestamp 1666464484
transform 1 0 25116 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_273
timestamp 1666464484
transform 1 0 26220 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_280
timestamp 1666464484
transform 1 0 26864 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_292
timestamp 1666464484
transform 1 0 27968 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_304
timestamp 1666464484
transform 1 0 29072 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_316
timestamp 1666464484
transform 1 0 30176 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_323
timestamp 1666464484
transform 1 0 30820 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_335
timestamp 1666464484
transform 1 0 31924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_347
timestamp 1666464484
transform 1 0 33028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_359
timestamp 1666464484
transform 1 0 34132 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_366
timestamp 1666464484
transform 1 0 34776 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_378
timestamp 1666464484
transform 1 0 35880 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_390
timestamp 1666464484
transform 1 0 36984 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_402
timestamp 1666464484
transform 1 0 38088 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_409
timestamp 1666464484
transform 1 0 38732 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1666464484
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1666464484
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_445
timestamp 1666464484
transform 1 0 42044 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_452
timestamp 1666464484
transform 1 0 42688 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_464
timestamp 1666464484
transform 1 0 43792 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_476
timestamp 1666464484
transform 1 0 44896 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_488
timestamp 1666464484
transform 1 0 46000 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_495
timestamp 1666464484
transform 1 0 46644 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_507
timestamp 1666464484
transform 1 0 47748 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_519
timestamp 1666464484
transform 1 0 48852 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_531
timestamp 1666464484
transform 1 0 49956 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_538
timestamp 1666464484
transform 1 0 50600 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_550
timestamp 1666464484
transform 1 0 51704 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_562
timestamp 1666464484
transform 1 0 52808 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_574
timestamp 1666464484
transform 1 0 53912 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_581
timestamp 1666464484
transform 1 0 54556 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_593
timestamp 1666464484
transform 1 0 55660 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_605
timestamp 1666464484
transform 1 0 56764 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_617
timestamp 1666464484
transform 1 0 57868 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_624
timestamp 1666464484
transform 1 0 58512 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1666464484
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1666464484
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1666464484
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_39
timestamp 1666464484
transform 1 0 4692 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_44
timestamp 1666464484
transform 1 0 5152 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_56
timestamp 1666464484
transform 1 0 6256 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_68
timestamp 1666464484
transform 1 0 7360 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_80
timestamp 1666464484
transform 1 0 8464 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_87
timestamp 1666464484
transform 1 0 9108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_99
timestamp 1666464484
transform 1 0 10212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_111
timestamp 1666464484
transform 1 0 11316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_123
timestamp 1666464484
transform 1 0 12420 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_130
timestamp 1666464484
transform 1 0 13064 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_142
timestamp 1666464484
transform 1 0 14168 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_154
timestamp 1666464484
transform 1 0 15272 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_166
timestamp 1666464484
transform 1 0 16376 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_173
timestamp 1666464484
transform 1 0 17020 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_185
timestamp 1666464484
transform 1 0 18124 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_197
timestamp 1666464484
transform 1 0 19228 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_209
timestamp 1666464484
transform 1 0 20332 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_216
timestamp 1666464484
transform 1 0 20976 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_228
timestamp 1666464484
transform 1 0 22080 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_240
timestamp 1666464484
transform 1 0 23184 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_252
timestamp 1666464484
transform 1 0 24288 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_259
timestamp 1666464484
transform 1 0 24932 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_271
timestamp 1666464484
transform 1 0 26036 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_283
timestamp 1666464484
transform 1 0 27140 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_295
timestamp 1666464484
transform 1 0 28244 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_302
timestamp 1666464484
transform 1 0 28888 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_314
timestamp 1666464484
transform 1 0 29992 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_326
timestamp 1666464484
transform 1 0 31096 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_338
timestamp 1666464484
transform 1 0 32200 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_345
timestamp 1666464484
transform 1 0 32844 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_357
timestamp 1666464484
transform 1 0 33948 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_369
timestamp 1666464484
transform 1 0 35052 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_381
timestamp 1666464484
transform 1 0 36156 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_388
timestamp 1666464484
transform 1 0 36800 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_400
timestamp 1666464484
transform 1 0 37904 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_412
timestamp 1666464484
transform 1 0 39008 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_424
timestamp 1666464484
transform 1 0 40112 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_431
timestamp 1666464484
transform 1 0 40756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_443
timestamp 1666464484
transform 1 0 41860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_455
timestamp 1666464484
transform 1 0 42964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_467
timestamp 1666464484
transform 1 0 44068 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_474
timestamp 1666464484
transform 1 0 44712 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_486
timestamp 1666464484
transform 1 0 45816 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_498
timestamp 1666464484
transform 1 0 46920 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_510
timestamp 1666464484
transform 1 0 48024 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1666464484
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1666464484
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1666464484
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1666464484
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_560
timestamp 1666464484
transform 1 0 52624 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_572
timestamp 1666464484
transform 1 0 53728 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_584
timestamp 1666464484
transform 1 0 54832 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_596
timestamp 1666464484
transform 1 0 55936 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_603
timestamp 1666464484
transform 1 0 56580 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_615
timestamp 1666464484
transform 1 0 57684 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_623
timestamp 1666464484
transform 1 0 58420 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1666464484
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_15
timestamp 1666464484
transform 1 0 2484 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_22
timestamp 1666464484
transform 1 0 3128 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_34
timestamp 1666464484
transform 1 0 4232 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_46
timestamp 1666464484
transform 1 0 5336 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_58
timestamp 1666464484
transform 1 0 6440 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1666464484
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_77
timestamp 1666464484
transform 1 0 8188 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_89
timestamp 1666464484
transform 1 0 9292 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_101
timestamp 1666464484
transform 1 0 10396 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_108
timestamp 1666464484
transform 1 0 11040 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_120
timestamp 1666464484
transform 1 0 12144 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_132
timestamp 1666464484
transform 1 0 13248 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_144
timestamp 1666464484
transform 1 0 14352 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_151
timestamp 1666464484
transform 1 0 14996 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_163
timestamp 1666464484
transform 1 0 16100 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_175
timestamp 1666464484
transform 1 0 17204 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_187
timestamp 1666464484
transform 1 0 18308 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_194
timestamp 1666464484
transform 1 0 18952 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_206
timestamp 1666464484
transform 1 0 20056 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_218
timestamp 1666464484
transform 1 0 21160 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_230
timestamp 1666464484
transform 1 0 22264 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_237
timestamp 1666464484
transform 1 0 22908 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_249
timestamp 1666464484
transform 1 0 24012 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_261
timestamp 1666464484
transform 1 0 25116 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_273
timestamp 1666464484
transform 1 0 26220 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_280
timestamp 1666464484
transform 1 0 26864 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_292
timestamp 1666464484
transform 1 0 27968 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_304
timestamp 1666464484
transform 1 0 29072 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_316
timestamp 1666464484
transform 1 0 30176 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_323
timestamp 1666464484
transform 1 0 30820 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_335
timestamp 1666464484
transform 1 0 31924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_347
timestamp 1666464484
transform 1 0 33028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_359
timestamp 1666464484
transform 1 0 34132 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_366
timestamp 1666464484
transform 1 0 34776 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_378
timestamp 1666464484
transform 1 0 35880 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_390
timestamp 1666464484
transform 1 0 36984 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_402
timestamp 1666464484
transform 1 0 38088 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_409
timestamp 1666464484
transform 1 0 38732 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1666464484
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1666464484
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_445
timestamp 1666464484
transform 1 0 42044 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_452
timestamp 1666464484
transform 1 0 42688 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_464
timestamp 1666464484
transform 1 0 43792 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_476
timestamp 1666464484
transform 1 0 44896 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_488
timestamp 1666464484
transform 1 0 46000 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_495
timestamp 1666464484
transform 1 0 46644 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_507
timestamp 1666464484
transform 1 0 47748 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_519
timestamp 1666464484
transform 1 0 48852 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_531
timestamp 1666464484
transform 1 0 49956 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_538
timestamp 1666464484
transform 1 0 50600 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_550
timestamp 1666464484
transform 1 0 51704 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_562
timestamp 1666464484
transform 1 0 52808 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_574
timestamp 1666464484
transform 1 0 53912 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_581
timestamp 1666464484
transform 1 0 54556 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_593
timestamp 1666464484
transform 1 0 55660 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_605
timestamp 1666464484
transform 1 0 56764 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_617
timestamp 1666464484
transform 1 0 57868 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_624
timestamp 1666464484
transform 1 0 58512 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1666464484
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1666464484
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1666464484
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_39
timestamp 1666464484
transform 1 0 4692 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_44
timestamp 1666464484
transform 1 0 5152 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_56
timestamp 1666464484
transform 1 0 6256 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_68
timestamp 1666464484
transform 1 0 7360 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_80
timestamp 1666464484
transform 1 0 8464 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_87
timestamp 1666464484
transform 1 0 9108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_99
timestamp 1666464484
transform 1 0 10212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_111
timestamp 1666464484
transform 1 0 11316 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_123
timestamp 1666464484
transform 1 0 12420 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_130
timestamp 1666464484
transform 1 0 13064 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_142
timestamp 1666464484
transform 1 0 14168 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_154
timestamp 1666464484
transform 1 0 15272 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_166
timestamp 1666464484
transform 1 0 16376 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_173
timestamp 1666464484
transform 1 0 17020 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_185
timestamp 1666464484
transform 1 0 18124 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_197
timestamp 1666464484
transform 1 0 19228 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_209
timestamp 1666464484
transform 1 0 20332 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_216
timestamp 1666464484
transform 1 0 20976 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_228
timestamp 1666464484
transform 1 0 22080 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_240
timestamp 1666464484
transform 1 0 23184 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_252
timestamp 1666464484
transform 1 0 24288 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_259
timestamp 1666464484
transform 1 0 24932 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_271
timestamp 1666464484
transform 1 0 26036 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_283
timestamp 1666464484
transform 1 0 27140 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_295
timestamp 1666464484
transform 1 0 28244 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_302
timestamp 1666464484
transform 1 0 28888 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_314
timestamp 1666464484
transform 1 0 29992 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_326
timestamp 1666464484
transform 1 0 31096 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_338
timestamp 1666464484
transform 1 0 32200 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_345
timestamp 1666464484
transform 1 0 32844 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_357
timestamp 1666464484
transform 1 0 33948 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_369
timestamp 1666464484
transform 1 0 35052 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_381
timestamp 1666464484
transform 1 0 36156 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_388
timestamp 1666464484
transform 1 0 36800 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_400
timestamp 1666464484
transform 1 0 37904 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_412
timestamp 1666464484
transform 1 0 39008 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_424
timestamp 1666464484
transform 1 0 40112 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_431
timestamp 1666464484
transform 1 0 40756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_443
timestamp 1666464484
transform 1 0 41860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_455
timestamp 1666464484
transform 1 0 42964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_467
timestamp 1666464484
transform 1 0 44068 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_474
timestamp 1666464484
transform 1 0 44712 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_486
timestamp 1666464484
transform 1 0 45816 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_498
timestamp 1666464484
transform 1 0 46920 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_510
timestamp 1666464484
transform 1 0 48024 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1666464484
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1666464484
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1666464484
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1666464484
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_560
timestamp 1666464484
transform 1 0 52624 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_572
timestamp 1666464484
transform 1 0 53728 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_584
timestamp 1666464484
transform 1 0 54832 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_596
timestamp 1666464484
transform 1 0 55936 0 -1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_603
timestamp 1666464484
transform 1 0 56580 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_615
timestamp 1666464484
transform 1 0 57684 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_623
timestamp 1666464484
transform 1 0 58420 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1666464484
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_15
timestamp 1666464484
transform 1 0 2484 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_22
timestamp 1666464484
transform 1 0 3128 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_34
timestamp 1666464484
transform 1 0 4232 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_46
timestamp 1666464484
transform 1 0 5336 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_58
timestamp 1666464484
transform 1 0 6440 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1666464484
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_77
timestamp 1666464484
transform 1 0 8188 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_89
timestamp 1666464484
transform 1 0 9292 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_101
timestamp 1666464484
transform 1 0 10396 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_108
timestamp 1666464484
transform 1 0 11040 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_120
timestamp 1666464484
transform 1 0 12144 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_132
timestamp 1666464484
transform 1 0 13248 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_144
timestamp 1666464484
transform 1 0 14352 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_151
timestamp 1666464484
transform 1 0 14996 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_163
timestamp 1666464484
transform 1 0 16100 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_175
timestamp 1666464484
transform 1 0 17204 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_187
timestamp 1666464484
transform 1 0 18308 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_194
timestamp 1666464484
transform 1 0 18952 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_206
timestamp 1666464484
transform 1 0 20056 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_218
timestamp 1666464484
transform 1 0 21160 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_230
timestamp 1666464484
transform 1 0 22264 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_237
timestamp 1666464484
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_249
timestamp 1666464484
transform 1 0 24012 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_261
timestamp 1666464484
transform 1 0 25116 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_273
timestamp 1666464484
transform 1 0 26220 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_280
timestamp 1666464484
transform 1 0 26864 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_292
timestamp 1666464484
transform 1 0 27968 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_304
timestamp 1666464484
transform 1 0 29072 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_316
timestamp 1666464484
transform 1 0 30176 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_323
timestamp 1666464484
transform 1 0 30820 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_335
timestamp 1666464484
transform 1 0 31924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_347
timestamp 1666464484
transform 1 0 33028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_359
timestamp 1666464484
transform 1 0 34132 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_366
timestamp 1666464484
transform 1 0 34776 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_378
timestamp 1666464484
transform 1 0 35880 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_390
timestamp 1666464484
transform 1 0 36984 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_402
timestamp 1666464484
transform 1 0 38088 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_409
timestamp 1666464484
transform 1 0 38732 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1666464484
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1666464484
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_445
timestamp 1666464484
transform 1 0 42044 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_452
timestamp 1666464484
transform 1 0 42688 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_464
timestamp 1666464484
transform 1 0 43792 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_476
timestamp 1666464484
transform 1 0 44896 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_488
timestamp 1666464484
transform 1 0 46000 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_495
timestamp 1666464484
transform 1 0 46644 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_507
timestamp 1666464484
transform 1 0 47748 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_519
timestamp 1666464484
transform 1 0 48852 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_531
timestamp 1666464484
transform 1 0 49956 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_538
timestamp 1666464484
transform 1 0 50600 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_550
timestamp 1666464484
transform 1 0 51704 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_562
timestamp 1666464484
transform 1 0 52808 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_574
timestamp 1666464484
transform 1 0 53912 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_581
timestamp 1666464484
transform 1 0 54556 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_593
timestamp 1666464484
transform 1 0 55660 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_605
timestamp 1666464484
transform 1 0 56764 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_617
timestamp 1666464484
transform 1 0 57868 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_624
timestamp 1666464484
transform 1 0 58512 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1666464484
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1666464484
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1666464484
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_39
timestamp 1666464484
transform 1 0 4692 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_44
timestamp 1666464484
transform 1 0 5152 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_56
timestamp 1666464484
transform 1 0 6256 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_68
timestamp 1666464484
transform 1 0 7360 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_80
timestamp 1666464484
transform 1 0 8464 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_87
timestamp 1666464484
transform 1 0 9108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_99
timestamp 1666464484
transform 1 0 10212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_111
timestamp 1666464484
transform 1 0 11316 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_123
timestamp 1666464484
transform 1 0 12420 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_130
timestamp 1666464484
transform 1 0 13064 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_142
timestamp 1666464484
transform 1 0 14168 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_154
timestamp 1666464484
transform 1 0 15272 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_166
timestamp 1666464484
transform 1 0 16376 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_173
timestamp 1666464484
transform 1 0 17020 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_185
timestamp 1666464484
transform 1 0 18124 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_197
timestamp 1666464484
transform 1 0 19228 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_209
timestamp 1666464484
transform 1 0 20332 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_216
timestamp 1666464484
transform 1 0 20976 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_228
timestamp 1666464484
transform 1 0 22080 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_240
timestamp 1666464484
transform 1 0 23184 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_252
timestamp 1666464484
transform 1 0 24288 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_259
timestamp 1666464484
transform 1 0 24932 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_271
timestamp 1666464484
transform 1 0 26036 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_283
timestamp 1666464484
transform 1 0 27140 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_295
timestamp 1666464484
transform 1 0 28244 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_302
timestamp 1666464484
transform 1 0 28888 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_314
timestamp 1666464484
transform 1 0 29992 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_326
timestamp 1666464484
transform 1 0 31096 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_338
timestamp 1666464484
transform 1 0 32200 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_345
timestamp 1666464484
transform 1 0 32844 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_357
timestamp 1666464484
transform 1 0 33948 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_369
timestamp 1666464484
transform 1 0 35052 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_381
timestamp 1666464484
transform 1 0 36156 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_388
timestamp 1666464484
transform 1 0 36800 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_400
timestamp 1666464484
transform 1 0 37904 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_412
timestamp 1666464484
transform 1 0 39008 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_424
timestamp 1666464484
transform 1 0 40112 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_431
timestamp 1666464484
transform 1 0 40756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_443
timestamp 1666464484
transform 1 0 41860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_455
timestamp 1666464484
transform 1 0 42964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_467
timestamp 1666464484
transform 1 0 44068 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_474
timestamp 1666464484
transform 1 0 44712 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_486
timestamp 1666464484
transform 1 0 45816 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_498
timestamp 1666464484
transform 1 0 46920 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_510
timestamp 1666464484
transform 1 0 48024 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1666464484
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1666464484
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1666464484
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1666464484
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_560
timestamp 1666464484
transform 1 0 52624 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_572
timestamp 1666464484
transform 1 0 53728 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_584
timestamp 1666464484
transform 1 0 54832 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_596
timestamp 1666464484
transform 1 0 55936 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_603
timestamp 1666464484
transform 1 0 56580 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_615
timestamp 1666464484
transform 1 0 57684 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_623
timestamp 1666464484
transform 1 0 58420 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1666464484
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_15
timestamp 1666464484
transform 1 0 2484 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_22
timestamp 1666464484
transform 1 0 3128 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_34
timestamp 1666464484
transform 1 0 4232 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_46
timestamp 1666464484
transform 1 0 5336 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_58
timestamp 1666464484
transform 1 0 6440 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1666464484
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_77
timestamp 1666464484
transform 1 0 8188 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_89
timestamp 1666464484
transform 1 0 9292 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_101
timestamp 1666464484
transform 1 0 10396 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_108
timestamp 1666464484
transform 1 0 11040 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_120
timestamp 1666464484
transform 1 0 12144 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_132
timestamp 1666464484
transform 1 0 13248 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_144
timestamp 1666464484
transform 1 0 14352 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_151
timestamp 1666464484
transform 1 0 14996 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_163
timestamp 1666464484
transform 1 0 16100 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_175
timestamp 1666464484
transform 1 0 17204 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_187
timestamp 1666464484
transform 1 0 18308 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_194
timestamp 1666464484
transform 1 0 18952 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_206
timestamp 1666464484
transform 1 0 20056 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_218
timestamp 1666464484
transform 1 0 21160 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_230
timestamp 1666464484
transform 1 0 22264 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_237
timestamp 1666464484
transform 1 0 22908 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_249
timestamp 1666464484
transform 1 0 24012 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_261
timestamp 1666464484
transform 1 0 25116 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_273
timestamp 1666464484
transform 1 0 26220 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_280
timestamp 1666464484
transform 1 0 26864 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_292
timestamp 1666464484
transform 1 0 27968 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_304
timestamp 1666464484
transform 1 0 29072 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_316
timestamp 1666464484
transform 1 0 30176 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_323
timestamp 1666464484
transform 1 0 30820 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_335
timestamp 1666464484
transform 1 0 31924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_347
timestamp 1666464484
transform 1 0 33028 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_359
timestamp 1666464484
transform 1 0 34132 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_366
timestamp 1666464484
transform 1 0 34776 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_378
timestamp 1666464484
transform 1 0 35880 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_390
timestamp 1666464484
transform 1 0 36984 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_402
timestamp 1666464484
transform 1 0 38088 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_409
timestamp 1666464484
transform 1 0 38732 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1666464484
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1666464484
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_445
timestamp 1666464484
transform 1 0 42044 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_452
timestamp 1666464484
transform 1 0 42688 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_464
timestamp 1666464484
transform 1 0 43792 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_476
timestamp 1666464484
transform 1 0 44896 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_488
timestamp 1666464484
transform 1 0 46000 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_495
timestamp 1666464484
transform 1 0 46644 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_507
timestamp 1666464484
transform 1 0 47748 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_519
timestamp 1666464484
transform 1 0 48852 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_531
timestamp 1666464484
transform 1 0 49956 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_538
timestamp 1666464484
transform 1 0 50600 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_550
timestamp 1666464484
transform 1 0 51704 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_562
timestamp 1666464484
transform 1 0 52808 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_574
timestamp 1666464484
transform 1 0 53912 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_581
timestamp 1666464484
transform 1 0 54556 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_593
timestamp 1666464484
transform 1 0 55660 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_605
timestamp 1666464484
transform 1 0 56764 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_617
timestamp 1666464484
transform 1 0 57868 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_624
timestamp 1666464484
transform 1 0 58512 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1666464484
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1666464484
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1666464484
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_39
timestamp 1666464484
transform 1 0 4692 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_44
timestamp 1666464484
transform 1 0 5152 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_56
timestamp 1666464484
transform 1 0 6256 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_68
timestamp 1666464484
transform 1 0 7360 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_80
timestamp 1666464484
transform 1 0 8464 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_87
timestamp 1666464484
transform 1 0 9108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_99
timestamp 1666464484
transform 1 0 10212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_111
timestamp 1666464484
transform 1 0 11316 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_123
timestamp 1666464484
transform 1 0 12420 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_130
timestamp 1666464484
transform 1 0 13064 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_142
timestamp 1666464484
transform 1 0 14168 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_154
timestamp 1666464484
transform 1 0 15272 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_166
timestamp 1666464484
transform 1 0 16376 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_173
timestamp 1666464484
transform 1 0 17020 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_185
timestamp 1666464484
transform 1 0 18124 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_197
timestamp 1666464484
transform 1 0 19228 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_209
timestamp 1666464484
transform 1 0 20332 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_216
timestamp 1666464484
transform 1 0 20976 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_228
timestamp 1666464484
transform 1 0 22080 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_240
timestamp 1666464484
transform 1 0 23184 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_252
timestamp 1666464484
transform 1 0 24288 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_259
timestamp 1666464484
transform 1 0 24932 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_271
timestamp 1666464484
transform 1 0 26036 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_283
timestamp 1666464484
transform 1 0 27140 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_295
timestamp 1666464484
transform 1 0 28244 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_302
timestamp 1666464484
transform 1 0 28888 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_314
timestamp 1666464484
transform 1 0 29992 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_326
timestamp 1666464484
transform 1 0 31096 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_338
timestamp 1666464484
transform 1 0 32200 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_345
timestamp 1666464484
transform 1 0 32844 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_357
timestamp 1666464484
transform 1 0 33948 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_369
timestamp 1666464484
transform 1 0 35052 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_381
timestamp 1666464484
transform 1 0 36156 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_388
timestamp 1666464484
transform 1 0 36800 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_400
timestamp 1666464484
transform 1 0 37904 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_412
timestamp 1666464484
transform 1 0 39008 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_424
timestamp 1666464484
transform 1 0 40112 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_431
timestamp 1666464484
transform 1 0 40756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_443
timestamp 1666464484
transform 1 0 41860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_455
timestamp 1666464484
transform 1 0 42964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_467
timestamp 1666464484
transform 1 0 44068 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_474
timestamp 1666464484
transform 1 0 44712 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_486
timestamp 1666464484
transform 1 0 45816 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_498
timestamp 1666464484
transform 1 0 46920 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_510
timestamp 1666464484
transform 1 0 48024 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1666464484
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1666464484
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1666464484
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1666464484
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_560
timestamp 1666464484
transform 1 0 52624 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_572
timestamp 1666464484
transform 1 0 53728 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_584
timestamp 1666464484
transform 1 0 54832 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_596
timestamp 1666464484
transform 1 0 55936 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_603
timestamp 1666464484
transform 1 0 56580 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_615
timestamp 1666464484
transform 1 0 57684 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_623
timestamp 1666464484
transform 1 0 58420 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1666464484
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_15
timestamp 1666464484
transform 1 0 2484 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_22
timestamp 1666464484
transform 1 0 3128 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_34
timestamp 1666464484
transform 1 0 4232 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_46
timestamp 1666464484
transform 1 0 5336 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_58
timestamp 1666464484
transform 1 0 6440 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1666464484
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_77
timestamp 1666464484
transform 1 0 8188 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_89
timestamp 1666464484
transform 1 0 9292 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_101
timestamp 1666464484
transform 1 0 10396 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_108
timestamp 1666464484
transform 1 0 11040 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_120
timestamp 1666464484
transform 1 0 12144 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_132
timestamp 1666464484
transform 1 0 13248 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_144
timestamp 1666464484
transform 1 0 14352 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_151
timestamp 1666464484
transform 1 0 14996 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_163
timestamp 1666464484
transform 1 0 16100 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_175
timestamp 1666464484
transform 1 0 17204 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_187
timestamp 1666464484
transform 1 0 18308 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_194
timestamp 1666464484
transform 1 0 18952 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_206
timestamp 1666464484
transform 1 0 20056 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_218
timestamp 1666464484
transform 1 0 21160 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_230
timestamp 1666464484
transform 1 0 22264 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_237
timestamp 1666464484
transform 1 0 22908 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_249
timestamp 1666464484
transform 1 0 24012 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_261
timestamp 1666464484
transform 1 0 25116 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_273
timestamp 1666464484
transform 1 0 26220 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_280
timestamp 1666464484
transform 1 0 26864 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_292
timestamp 1666464484
transform 1 0 27968 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_304
timestamp 1666464484
transform 1 0 29072 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_316
timestamp 1666464484
transform 1 0 30176 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_323
timestamp 1666464484
transform 1 0 30820 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_335
timestamp 1666464484
transform 1 0 31924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_347
timestamp 1666464484
transform 1 0 33028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_359
timestamp 1666464484
transform 1 0 34132 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_366
timestamp 1666464484
transform 1 0 34776 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_378
timestamp 1666464484
transform 1 0 35880 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_390
timestamp 1666464484
transform 1 0 36984 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_402
timestamp 1666464484
transform 1 0 38088 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_409
timestamp 1666464484
transform 1 0 38732 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1666464484
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1666464484
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_445
timestamp 1666464484
transform 1 0 42044 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_452
timestamp 1666464484
transform 1 0 42688 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_464
timestamp 1666464484
transform 1 0 43792 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_476
timestamp 1666464484
transform 1 0 44896 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_488
timestamp 1666464484
transform 1 0 46000 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_495
timestamp 1666464484
transform 1 0 46644 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_507
timestamp 1666464484
transform 1 0 47748 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_519
timestamp 1666464484
transform 1 0 48852 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_531
timestamp 1666464484
transform 1 0 49956 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_538
timestamp 1666464484
transform 1 0 50600 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_550
timestamp 1666464484
transform 1 0 51704 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_562
timestamp 1666464484
transform 1 0 52808 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_574
timestamp 1666464484
transform 1 0 53912 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_581
timestamp 1666464484
transform 1 0 54556 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_593
timestamp 1666464484
transform 1 0 55660 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_605
timestamp 1666464484
transform 1 0 56764 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_617
timestamp 1666464484
transform 1 0 57868 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_624
timestamp 1666464484
transform 1 0 58512 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1666464484
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1666464484
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1666464484
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_39
timestamp 1666464484
transform 1 0 4692 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_44
timestamp 1666464484
transform 1 0 5152 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_56
timestamp 1666464484
transform 1 0 6256 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_68
timestamp 1666464484
transform 1 0 7360 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_80
timestamp 1666464484
transform 1 0 8464 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_87
timestamp 1666464484
transform 1 0 9108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_99
timestamp 1666464484
transform 1 0 10212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_111
timestamp 1666464484
transform 1 0 11316 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_123
timestamp 1666464484
transform 1 0 12420 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_130
timestamp 1666464484
transform 1 0 13064 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_142
timestamp 1666464484
transform 1 0 14168 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_154
timestamp 1666464484
transform 1 0 15272 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_166
timestamp 1666464484
transform 1 0 16376 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_173
timestamp 1666464484
transform 1 0 17020 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_185
timestamp 1666464484
transform 1 0 18124 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_197
timestamp 1666464484
transform 1 0 19228 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_209
timestamp 1666464484
transform 1 0 20332 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_216
timestamp 1666464484
transform 1 0 20976 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_228
timestamp 1666464484
transform 1 0 22080 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_240
timestamp 1666464484
transform 1 0 23184 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_252
timestamp 1666464484
transform 1 0 24288 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_259
timestamp 1666464484
transform 1 0 24932 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_271
timestamp 1666464484
transform 1 0 26036 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_283
timestamp 1666464484
transform 1 0 27140 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_295
timestamp 1666464484
transform 1 0 28244 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_302
timestamp 1666464484
transform 1 0 28888 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_314
timestamp 1666464484
transform 1 0 29992 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_326
timestamp 1666464484
transform 1 0 31096 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_338
timestamp 1666464484
transform 1 0 32200 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_345
timestamp 1666464484
transform 1 0 32844 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_357
timestamp 1666464484
transform 1 0 33948 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_369
timestamp 1666464484
transform 1 0 35052 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_381
timestamp 1666464484
transform 1 0 36156 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_388
timestamp 1666464484
transform 1 0 36800 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_400
timestamp 1666464484
transform 1 0 37904 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_412
timestamp 1666464484
transform 1 0 39008 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_424
timestamp 1666464484
transform 1 0 40112 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_431
timestamp 1666464484
transform 1 0 40756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_443
timestamp 1666464484
transform 1 0 41860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_455
timestamp 1666464484
transform 1 0 42964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_467
timestamp 1666464484
transform 1 0 44068 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_474
timestamp 1666464484
transform 1 0 44712 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_486
timestamp 1666464484
transform 1 0 45816 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_498
timestamp 1666464484
transform 1 0 46920 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_510
timestamp 1666464484
transform 1 0 48024 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1666464484
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1666464484
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1666464484
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1666464484
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_560
timestamp 1666464484
transform 1 0 52624 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_572
timestamp 1666464484
transform 1 0 53728 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_584
timestamp 1666464484
transform 1 0 54832 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_596
timestamp 1666464484
transform 1 0 55936 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_603
timestamp 1666464484
transform 1 0 56580 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_615
timestamp 1666464484
transform 1 0 57684 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_623
timestamp 1666464484
transform 1 0 58420 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1666464484
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_15
timestamp 1666464484
transform 1 0 2484 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_22
timestamp 1666464484
transform 1 0 3128 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_34
timestamp 1666464484
transform 1 0 4232 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_46
timestamp 1666464484
transform 1 0 5336 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_58
timestamp 1666464484
transform 1 0 6440 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1666464484
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_77
timestamp 1666464484
transform 1 0 8188 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_89
timestamp 1666464484
transform 1 0 9292 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_101
timestamp 1666464484
transform 1 0 10396 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_108
timestamp 1666464484
transform 1 0 11040 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_120
timestamp 1666464484
transform 1 0 12144 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_132
timestamp 1666464484
transform 1 0 13248 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_144
timestamp 1666464484
transform 1 0 14352 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_151
timestamp 1666464484
transform 1 0 14996 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_163
timestamp 1666464484
transform 1 0 16100 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_175
timestamp 1666464484
transform 1 0 17204 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_187
timestamp 1666464484
transform 1 0 18308 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_194
timestamp 1666464484
transform 1 0 18952 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_206
timestamp 1666464484
transform 1 0 20056 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_218
timestamp 1666464484
transform 1 0 21160 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_230
timestamp 1666464484
transform 1 0 22264 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_237
timestamp 1666464484
transform 1 0 22908 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_249
timestamp 1666464484
transform 1 0 24012 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_261
timestamp 1666464484
transform 1 0 25116 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_273
timestamp 1666464484
transform 1 0 26220 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_280
timestamp 1666464484
transform 1 0 26864 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_292
timestamp 1666464484
transform 1 0 27968 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_304
timestamp 1666464484
transform 1 0 29072 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_316
timestamp 1666464484
transform 1 0 30176 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_323
timestamp 1666464484
transform 1 0 30820 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_335
timestamp 1666464484
transform 1 0 31924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_347
timestamp 1666464484
transform 1 0 33028 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_359
timestamp 1666464484
transform 1 0 34132 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_366
timestamp 1666464484
transform 1 0 34776 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_378
timestamp 1666464484
transform 1 0 35880 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_390
timestamp 1666464484
transform 1 0 36984 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_402
timestamp 1666464484
transform 1 0 38088 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_409
timestamp 1666464484
transform 1 0 38732 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1666464484
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1666464484
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_445
timestamp 1666464484
transform 1 0 42044 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_452
timestamp 1666464484
transform 1 0 42688 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_464
timestamp 1666464484
transform 1 0 43792 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_476
timestamp 1666464484
transform 1 0 44896 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_488
timestamp 1666464484
transform 1 0 46000 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_495
timestamp 1666464484
transform 1 0 46644 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_507
timestamp 1666464484
transform 1 0 47748 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_519
timestamp 1666464484
transform 1 0 48852 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_531
timestamp 1666464484
transform 1 0 49956 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_538
timestamp 1666464484
transform 1 0 50600 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_550
timestamp 1666464484
transform 1 0 51704 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_562
timestamp 1666464484
transform 1 0 52808 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_574
timestamp 1666464484
transform 1 0 53912 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_581
timestamp 1666464484
transform 1 0 54556 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_593
timestamp 1666464484
transform 1 0 55660 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_605
timestamp 1666464484
transform 1 0 56764 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_617
timestamp 1666464484
transform 1 0 57868 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_624
timestamp 1666464484
transform 1 0 58512 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1666464484
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1666464484
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1666464484
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_39
timestamp 1666464484
transform 1 0 4692 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_44
timestamp 1666464484
transform 1 0 5152 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_56
timestamp 1666464484
transform 1 0 6256 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_68
timestamp 1666464484
transform 1 0 7360 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_80
timestamp 1666464484
transform 1 0 8464 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_87
timestamp 1666464484
transform 1 0 9108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_99
timestamp 1666464484
transform 1 0 10212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_111
timestamp 1666464484
transform 1 0 11316 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_123
timestamp 1666464484
transform 1 0 12420 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_130
timestamp 1666464484
transform 1 0 13064 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_142
timestamp 1666464484
transform 1 0 14168 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_154
timestamp 1666464484
transform 1 0 15272 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_166
timestamp 1666464484
transform 1 0 16376 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_173
timestamp 1666464484
transform 1 0 17020 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_185
timestamp 1666464484
transform 1 0 18124 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_197
timestamp 1666464484
transform 1 0 19228 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_209
timestamp 1666464484
transform 1 0 20332 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_216
timestamp 1666464484
transform 1 0 20976 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_228
timestamp 1666464484
transform 1 0 22080 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_240
timestamp 1666464484
transform 1 0 23184 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_252
timestamp 1666464484
transform 1 0 24288 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_259
timestamp 1666464484
transform 1 0 24932 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_271
timestamp 1666464484
transform 1 0 26036 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_283
timestamp 1666464484
transform 1 0 27140 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_295
timestamp 1666464484
transform 1 0 28244 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_302
timestamp 1666464484
transform 1 0 28888 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_314
timestamp 1666464484
transform 1 0 29992 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_326
timestamp 1666464484
transform 1 0 31096 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_338
timestamp 1666464484
transform 1 0 32200 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_345
timestamp 1666464484
transform 1 0 32844 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_357
timestamp 1666464484
transform 1 0 33948 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_369
timestamp 1666464484
transform 1 0 35052 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_381
timestamp 1666464484
transform 1 0 36156 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_388
timestamp 1666464484
transform 1 0 36800 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_400
timestamp 1666464484
transform 1 0 37904 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_412
timestamp 1666464484
transform 1 0 39008 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_424
timestamp 1666464484
transform 1 0 40112 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_431
timestamp 1666464484
transform 1 0 40756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_443
timestamp 1666464484
transform 1 0 41860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_455
timestamp 1666464484
transform 1 0 42964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_467
timestamp 1666464484
transform 1 0 44068 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_474
timestamp 1666464484
transform 1 0 44712 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_486
timestamp 1666464484
transform 1 0 45816 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_498
timestamp 1666464484
transform 1 0 46920 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_510
timestamp 1666464484
transform 1 0 48024 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1666464484
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1666464484
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1666464484
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1666464484
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_560
timestamp 1666464484
transform 1 0 52624 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_572
timestamp 1666464484
transform 1 0 53728 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_584
timestamp 1666464484
transform 1 0 54832 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_596
timestamp 1666464484
transform 1 0 55936 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_603
timestamp 1666464484
transform 1 0 56580 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_615
timestamp 1666464484
transform 1 0 57684 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_623
timestamp 1666464484
transform 1 0 58420 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1666464484
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_15
timestamp 1666464484
transform 1 0 2484 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_22
timestamp 1666464484
transform 1 0 3128 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_34
timestamp 1666464484
transform 1 0 4232 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_46
timestamp 1666464484
transform 1 0 5336 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_58
timestamp 1666464484
transform 1 0 6440 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1666464484
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_77
timestamp 1666464484
transform 1 0 8188 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_89
timestamp 1666464484
transform 1 0 9292 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_101
timestamp 1666464484
transform 1 0 10396 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_108
timestamp 1666464484
transform 1 0 11040 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_120
timestamp 1666464484
transform 1 0 12144 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_132
timestamp 1666464484
transform 1 0 13248 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_144
timestamp 1666464484
transform 1 0 14352 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_151
timestamp 1666464484
transform 1 0 14996 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_163
timestamp 1666464484
transform 1 0 16100 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_175
timestamp 1666464484
transform 1 0 17204 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_187
timestamp 1666464484
transform 1 0 18308 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_194
timestamp 1666464484
transform 1 0 18952 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_206
timestamp 1666464484
transform 1 0 20056 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_218
timestamp 1666464484
transform 1 0 21160 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_230
timestamp 1666464484
transform 1 0 22264 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_237
timestamp 1666464484
transform 1 0 22908 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_249
timestamp 1666464484
transform 1 0 24012 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_261
timestamp 1666464484
transform 1 0 25116 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_273
timestamp 1666464484
transform 1 0 26220 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_280
timestamp 1666464484
transform 1 0 26864 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_292
timestamp 1666464484
transform 1 0 27968 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_304
timestamp 1666464484
transform 1 0 29072 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_316
timestamp 1666464484
transform 1 0 30176 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_323
timestamp 1666464484
transform 1 0 30820 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_335
timestamp 1666464484
transform 1 0 31924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_347
timestamp 1666464484
transform 1 0 33028 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_359
timestamp 1666464484
transform 1 0 34132 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_366
timestamp 1666464484
transform 1 0 34776 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_378
timestamp 1666464484
transform 1 0 35880 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_390
timestamp 1666464484
transform 1 0 36984 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_402
timestamp 1666464484
transform 1 0 38088 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_409
timestamp 1666464484
transform 1 0 38732 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1666464484
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1666464484
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_445
timestamp 1666464484
transform 1 0 42044 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_452
timestamp 1666464484
transform 1 0 42688 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_464
timestamp 1666464484
transform 1 0 43792 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_476
timestamp 1666464484
transform 1 0 44896 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_488
timestamp 1666464484
transform 1 0 46000 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_495
timestamp 1666464484
transform 1 0 46644 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_507
timestamp 1666464484
transform 1 0 47748 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_519
timestamp 1666464484
transform 1 0 48852 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_531
timestamp 1666464484
transform 1 0 49956 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_538
timestamp 1666464484
transform 1 0 50600 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_550
timestamp 1666464484
transform 1 0 51704 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_562
timestamp 1666464484
transform 1 0 52808 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_574
timestamp 1666464484
transform 1 0 53912 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_581
timestamp 1666464484
transform 1 0 54556 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_593
timestamp 1666464484
transform 1 0 55660 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_605
timestamp 1666464484
transform 1 0 56764 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_617
timestamp 1666464484
transform 1 0 57868 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_624
timestamp 1666464484
transform 1 0 58512 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1666464484
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1666464484
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1666464484
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_39
timestamp 1666464484
transform 1 0 4692 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_44
timestamp 1666464484
transform 1 0 5152 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_56
timestamp 1666464484
transform 1 0 6256 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_68
timestamp 1666464484
transform 1 0 7360 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_80
timestamp 1666464484
transform 1 0 8464 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_87
timestamp 1666464484
transform 1 0 9108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_99
timestamp 1666464484
transform 1 0 10212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_111
timestamp 1666464484
transform 1 0 11316 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_123
timestamp 1666464484
transform 1 0 12420 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_130
timestamp 1666464484
transform 1 0 13064 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_142
timestamp 1666464484
transform 1 0 14168 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_154
timestamp 1666464484
transform 1 0 15272 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_166
timestamp 1666464484
transform 1 0 16376 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_173
timestamp 1666464484
transform 1 0 17020 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_185
timestamp 1666464484
transform 1 0 18124 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_197
timestamp 1666464484
transform 1 0 19228 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_209
timestamp 1666464484
transform 1 0 20332 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_216
timestamp 1666464484
transform 1 0 20976 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_228
timestamp 1666464484
transform 1 0 22080 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_240
timestamp 1666464484
transform 1 0 23184 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_252
timestamp 1666464484
transform 1 0 24288 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_259
timestamp 1666464484
transform 1 0 24932 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_271
timestamp 1666464484
transform 1 0 26036 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_283
timestamp 1666464484
transform 1 0 27140 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_295
timestamp 1666464484
transform 1 0 28244 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_302
timestamp 1666464484
transform 1 0 28888 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_314
timestamp 1666464484
transform 1 0 29992 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_326
timestamp 1666464484
transform 1 0 31096 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_338
timestamp 1666464484
transform 1 0 32200 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_345
timestamp 1666464484
transform 1 0 32844 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_357
timestamp 1666464484
transform 1 0 33948 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_369
timestamp 1666464484
transform 1 0 35052 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_381
timestamp 1666464484
transform 1 0 36156 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_388
timestamp 1666464484
transform 1 0 36800 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_400
timestamp 1666464484
transform 1 0 37904 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_412
timestamp 1666464484
transform 1 0 39008 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_424
timestamp 1666464484
transform 1 0 40112 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_431
timestamp 1666464484
transform 1 0 40756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_443
timestamp 1666464484
transform 1 0 41860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_455
timestamp 1666464484
transform 1 0 42964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_467
timestamp 1666464484
transform 1 0 44068 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_474
timestamp 1666464484
transform 1 0 44712 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_486
timestamp 1666464484
transform 1 0 45816 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_498
timestamp 1666464484
transform 1 0 46920 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_510
timestamp 1666464484
transform 1 0 48024 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1666464484
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1666464484
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1666464484
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1666464484
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_560
timestamp 1666464484
transform 1 0 52624 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_572
timestamp 1666464484
transform 1 0 53728 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_584
timestamp 1666464484
transform 1 0 54832 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_596
timestamp 1666464484
transform 1 0 55936 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_603
timestamp 1666464484
transform 1 0 56580 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_615
timestamp 1666464484
transform 1 0 57684 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_623
timestamp 1666464484
transform 1 0 58420 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1666464484
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_15
timestamp 1666464484
transform 1 0 2484 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_22
timestamp 1666464484
transform 1 0 3128 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_34
timestamp 1666464484
transform 1 0 4232 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_46
timestamp 1666464484
transform 1 0 5336 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_58
timestamp 1666464484
transform 1 0 6440 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1666464484
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_77
timestamp 1666464484
transform 1 0 8188 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_89
timestamp 1666464484
transform 1 0 9292 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_101
timestamp 1666464484
transform 1 0 10396 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_108
timestamp 1666464484
transform 1 0 11040 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_120
timestamp 1666464484
transform 1 0 12144 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_132
timestamp 1666464484
transform 1 0 13248 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_144
timestamp 1666464484
transform 1 0 14352 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_151
timestamp 1666464484
transform 1 0 14996 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_163
timestamp 1666464484
transform 1 0 16100 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_175
timestamp 1666464484
transform 1 0 17204 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_187
timestamp 1666464484
transform 1 0 18308 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_194
timestamp 1666464484
transform 1 0 18952 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_206
timestamp 1666464484
transform 1 0 20056 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_218
timestamp 1666464484
transform 1 0 21160 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_230
timestamp 1666464484
transform 1 0 22264 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_237
timestamp 1666464484
transform 1 0 22908 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_249
timestamp 1666464484
transform 1 0 24012 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_261
timestamp 1666464484
transform 1 0 25116 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_273
timestamp 1666464484
transform 1 0 26220 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_280
timestamp 1666464484
transform 1 0 26864 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_292
timestamp 1666464484
transform 1 0 27968 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_304
timestamp 1666464484
transform 1 0 29072 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_308
timestamp 1666464484
transform 1 0 29440 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_320
timestamp 1666464484
transform 1 0 30544 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_323
timestamp 1666464484
transform 1 0 30820 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_335
timestamp 1666464484
transform 1 0 31924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_347
timestamp 1666464484
transform 1 0 33028 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_359
timestamp 1666464484
transform 1 0 34132 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_92_366
timestamp 1666464484
transform 1 0 34776 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_92_370
timestamp 1666464484
transform 1 0 35144 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_378
timestamp 1666464484
transform 1 0 35880 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_381
timestamp 1666464484
transform 1 0 36156 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_393
timestamp 1666464484
transform 1 0 37260 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_405
timestamp 1666464484
transform 1 0 38364 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_409
timestamp 1666464484
transform 1 0 38732 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1666464484
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1666464484
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_445
timestamp 1666464484
transform 1 0 42044 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_452
timestamp 1666464484
transform 1 0 42688 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_464
timestamp 1666464484
transform 1 0 43792 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_476
timestamp 1666464484
transform 1 0 44896 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_488
timestamp 1666464484
transform 1 0 46000 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_495
timestamp 1666464484
transform 1 0 46644 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_507
timestamp 1666464484
transform 1 0 47748 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_519
timestamp 1666464484
transform 1 0 48852 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_531
timestamp 1666464484
transform 1 0 49956 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_538
timestamp 1666464484
transform 1 0 50600 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_550
timestamp 1666464484
transform 1 0 51704 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_562
timestamp 1666464484
transform 1 0 52808 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_574
timestamp 1666464484
transform 1 0 53912 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_581
timestamp 1666464484
transform 1 0 54556 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_593
timestamp 1666464484
transform 1 0 55660 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_605
timestamp 1666464484
transform 1 0 56764 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_617
timestamp 1666464484
transform 1 0 57868 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_624
timestamp 1666464484
transform 1 0 58512 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1666464484
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1666464484
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1666464484
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_39
timestamp 1666464484
transform 1 0 4692 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_44
timestamp 1666464484
transform 1 0 5152 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_56
timestamp 1666464484
transform 1 0 6256 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_68
timestamp 1666464484
transform 1 0 7360 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_80
timestamp 1666464484
transform 1 0 8464 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_87
timestamp 1666464484
transform 1 0 9108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_99
timestamp 1666464484
transform 1 0 10212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_111
timestamp 1666464484
transform 1 0 11316 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_123
timestamp 1666464484
transform 1 0 12420 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_130
timestamp 1666464484
transform 1 0 13064 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_142
timestamp 1666464484
transform 1 0 14168 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_154
timestamp 1666464484
transform 1 0 15272 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_166
timestamp 1666464484
transform 1 0 16376 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_173
timestamp 1666464484
transform 1 0 17020 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_185
timestamp 1666464484
transform 1 0 18124 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_197
timestamp 1666464484
transform 1 0 19228 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_209
timestamp 1666464484
transform 1 0 20332 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_216
timestamp 1666464484
transform 1 0 20976 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_228
timestamp 1666464484
transform 1 0 22080 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_240
timestamp 1666464484
transform 1 0 23184 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_252
timestamp 1666464484
transform 1 0 24288 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_259
timestamp 1666464484
transform 1 0 24932 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_271
timestamp 1666464484
transform 1 0 26036 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_283
timestamp 1666464484
transform 1 0 27140 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_295
timestamp 1666464484
transform 1 0 28244 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_93_302
timestamp 1666464484
transform 1 0 28888 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_308
timestamp 1666464484
transform 1 0 29440 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_312
timestamp 1666464484
transform 1 0 29808 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_318
timestamp 1666464484
transform 1 0 30360 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_330
timestamp 1666464484
transform 1 0 31464 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_342
timestamp 1666464484
transform 1 0 32568 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_345
timestamp 1666464484
transform 1 0 32844 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_349
timestamp 1666464484
transform 1 0 33212 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_355
timestamp 1666464484
transform 1 0 33764 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_359
timestamp 1666464484
transform 1 0 34132 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_93_381
timestamp 1666464484
transform 1 0 36156 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_388
timestamp 1666464484
transform 1 0 36800 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_400
timestamp 1666464484
transform 1 0 37904 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_408
timestamp 1666464484
transform 1 0 38640 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_93_414
timestamp 1666464484
transform 1 0 39192 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_420
timestamp 1666464484
transform 1 0 39744 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_93_423
timestamp 1666464484
transform 1 0 40020 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_429
timestamp 1666464484
transform 1 0 40572 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_431
timestamp 1666464484
transform 1 0 40756 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_435
timestamp 1666464484
transform 1 0 41124 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_447
timestamp 1666464484
transform 1 0 42228 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_459
timestamp 1666464484
transform 1 0 43332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_471
timestamp 1666464484
transform 1 0 44436 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_474
timestamp 1666464484
transform 1 0 44712 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_486
timestamp 1666464484
transform 1 0 45816 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_498
timestamp 1666464484
transform 1 0 46920 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_510
timestamp 1666464484
transform 1 0 48024 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1666464484
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1666464484
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1666464484
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1666464484
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_560
timestamp 1666464484
transform 1 0 52624 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_572
timestamp 1666464484
transform 1 0 53728 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_584
timestamp 1666464484
transform 1 0 54832 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_596
timestamp 1666464484
transform 1 0 55936 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_603
timestamp 1666464484
transform 1 0 56580 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_615
timestamp 1666464484
transform 1 0 57684 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_623
timestamp 1666464484
transform 1 0 58420 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1666464484
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_15
timestamp 1666464484
transform 1 0 2484 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_22
timestamp 1666464484
transform 1 0 3128 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_34
timestamp 1666464484
transform 1 0 4232 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_46
timestamp 1666464484
transform 1 0 5336 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_58
timestamp 1666464484
transform 1 0 6440 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1666464484
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_77
timestamp 1666464484
transform 1 0 8188 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_89
timestamp 1666464484
transform 1 0 9292 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_101
timestamp 1666464484
transform 1 0 10396 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_108
timestamp 1666464484
transform 1 0 11040 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_120
timestamp 1666464484
transform 1 0 12144 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_132
timestamp 1666464484
transform 1 0 13248 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_144
timestamp 1666464484
transform 1 0 14352 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_151
timestamp 1666464484
transform 1 0 14996 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_163
timestamp 1666464484
transform 1 0 16100 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_175
timestamp 1666464484
transform 1 0 17204 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_187
timestamp 1666464484
transform 1 0 18308 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_194
timestamp 1666464484
transform 1 0 18952 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_206
timestamp 1666464484
transform 1 0 20056 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_218
timestamp 1666464484
transform 1 0 21160 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_230
timestamp 1666464484
transform 1 0 22264 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_237
timestamp 1666464484
transform 1 0 22908 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_249
timestamp 1666464484
transform 1 0 24012 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_261
timestamp 1666464484
transform 1 0 25116 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_273
timestamp 1666464484
transform 1 0 26220 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_280
timestamp 1666464484
transform 1 0 26864 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_94_292
timestamp 1666464484
transform 1 0 27968 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_296
timestamp 1666464484
transform 1 0 28336 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_302
timestamp 1666464484
transform 1 0 28888 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_309
timestamp 1666464484
transform 1 0 29532 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_313
timestamp 1666464484
transform 1 0 29900 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_317
timestamp 1666464484
transform 1 0 30268 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_321
timestamp 1666464484
transform 1 0 30636 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_323
timestamp 1666464484
transform 1 0 30820 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_327
timestamp 1666464484
transform 1 0 31188 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_330
timestamp 1666464484
transform 1 0 31464 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_336
timestamp 1666464484
transform 1 0 32016 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_342
timestamp 1666464484
transform 1 0 32568 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_349
timestamp 1666464484
transform 1 0 33212 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_358
timestamp 1666464484
transform 1 0 34040 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_364
timestamp 1666464484
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_366
timestamp 1666464484
transform 1 0 34776 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_371
timestamp 1666464484
transform 1 0 35236 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_375
timestamp 1666464484
transform 1 0 35604 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_378
timestamp 1666464484
transform 1 0 35880 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_384
timestamp 1666464484
transform 1 0 36432 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_390
timestamp 1666464484
transform 1 0 36984 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_398
timestamp 1666464484
transform 1 0 37720 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_402
timestamp 1666464484
transform 1 0 38088 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_94_409
timestamp 1666464484
transform 1 0 38732 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_414
timestamp 1666464484
transform 1 0 39192 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_421
timestamp 1666464484
transform 1 0 39836 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_427
timestamp 1666464484
transform 1 0 40388 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_433
timestamp 1666464484
transform 1 0 40940 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_439
timestamp 1666464484
transform 1 0 41492 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_452
timestamp 1666464484
transform 1 0 42688 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_464
timestamp 1666464484
transform 1 0 43792 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_476
timestamp 1666464484
transform 1 0 44896 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_488
timestamp 1666464484
transform 1 0 46000 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_495
timestamp 1666464484
transform 1 0 46644 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_507
timestamp 1666464484
transform 1 0 47748 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_519
timestamp 1666464484
transform 1 0 48852 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_531
timestamp 1666464484
transform 1 0 49956 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_538
timestamp 1666464484
transform 1 0 50600 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_550
timestamp 1666464484
transform 1 0 51704 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_562
timestamp 1666464484
transform 1 0 52808 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_574
timestamp 1666464484
transform 1 0 53912 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_581
timestamp 1666464484
transform 1 0 54556 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_593
timestamp 1666464484
transform 1 0 55660 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_605
timestamp 1666464484
transform 1 0 56764 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_617
timestamp 1666464484
transform 1 0 57868 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_624
timestamp 1666464484
transform 1 0 58512 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1666464484
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1666464484
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1666464484
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_39
timestamp 1666464484
transform 1 0 4692 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_44
timestamp 1666464484
transform 1 0 5152 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_56
timestamp 1666464484
transform 1 0 6256 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_68
timestamp 1666464484
transform 1 0 7360 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_80
timestamp 1666464484
transform 1 0 8464 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_87
timestamp 1666464484
transform 1 0 9108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_99
timestamp 1666464484
transform 1 0 10212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_111
timestamp 1666464484
transform 1 0 11316 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_123
timestamp 1666464484
transform 1 0 12420 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_130
timestamp 1666464484
transform 1 0 13064 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_142
timestamp 1666464484
transform 1 0 14168 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_154
timestamp 1666464484
transform 1 0 15272 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_166
timestamp 1666464484
transform 1 0 16376 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_173
timestamp 1666464484
transform 1 0 17020 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_185
timestamp 1666464484
transform 1 0 18124 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_197
timestamp 1666464484
transform 1 0 19228 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_209
timestamp 1666464484
transform 1 0 20332 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_216
timestamp 1666464484
transform 1 0 20976 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_228
timestamp 1666464484
transform 1 0 22080 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_240
timestamp 1666464484
transform 1 0 23184 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_252
timestamp 1666464484
transform 1 0 24288 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_95_259
timestamp 1666464484
transform 1 0 24932 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_267
timestamp 1666464484
transform 1 0 25668 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_271
timestamp 1666464484
transform 1 0 26036 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_277
timestamp 1666464484
transform 1 0 26588 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_283
timestamp 1666464484
transform 1 0 27140 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_286
timestamp 1666464484
transform 1 0 27416 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_292
timestamp 1666464484
transform 1 0 27968 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_299
timestamp 1666464484
transform 1 0 28612 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_302
timestamp 1666464484
transform 1 0 28888 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_306
timestamp 1666464484
transform 1 0 29256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_311
timestamp 1666464484
transform 1 0 29716 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_320
timestamp 1666464484
transform 1 0 30544 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_328
timestamp 1666464484
transform 1 0 31280 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_342
timestamp 1666464484
transform 1 0 32568 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_345
timestamp 1666464484
transform 1 0 32844 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_351
timestamp 1666464484
transform 1 0 33396 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_359
timestamp 1666464484
transform 1 0 34132 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_369
timestamp 1666464484
transform 1 0 35052 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_376
timestamp 1666464484
transform 1 0 35696 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_383
timestamp 1666464484
transform 1 0 36340 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_388
timestamp 1666464484
transform 1 0 36800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_393
timestamp 1666464484
transform 1 0 37260 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_399
timestamp 1666464484
transform 1 0 37812 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_408
timestamp 1666464484
transform 1 0 38640 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_416
timestamp 1666464484
transform 1 0 39376 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_421
timestamp 1666464484
transform 1 0 39836 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_428
timestamp 1666464484
transform 1 0 40480 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_431
timestamp 1666464484
transform 1 0 40756 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_436
timestamp 1666464484
transform 1 0 41216 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_448
timestamp 1666464484
transform 1 0 42320 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_454
timestamp 1666464484
transform 1 0 42872 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_466
timestamp 1666464484
transform 1 0 43976 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_472
timestamp 1666464484
transform 1 0 44528 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_474
timestamp 1666464484
transform 1 0 44712 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_486
timestamp 1666464484
transform 1 0 45816 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_498
timestamp 1666464484
transform 1 0 46920 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_510
timestamp 1666464484
transform 1 0 48024 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1666464484
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1666464484
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1666464484
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1666464484
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_560
timestamp 1666464484
transform 1 0 52624 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_572
timestamp 1666464484
transform 1 0 53728 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_584
timestamp 1666464484
transform 1 0 54832 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_596
timestamp 1666464484
transform 1 0 55936 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_603
timestamp 1666464484
transform 1 0 56580 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_615
timestamp 1666464484
transform 1 0 57684 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_623
timestamp 1666464484
transform 1 0 58420 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1666464484
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_15
timestamp 1666464484
transform 1 0 2484 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_22
timestamp 1666464484
transform 1 0 3128 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_34
timestamp 1666464484
transform 1 0 4232 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_46
timestamp 1666464484
transform 1 0 5336 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_58
timestamp 1666464484
transform 1 0 6440 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1666464484
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_77
timestamp 1666464484
transform 1 0 8188 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_89
timestamp 1666464484
transform 1 0 9292 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_101
timestamp 1666464484
transform 1 0 10396 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_108
timestamp 1666464484
transform 1 0 11040 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_120
timestamp 1666464484
transform 1 0 12144 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_132
timestamp 1666464484
transform 1 0 13248 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_144
timestamp 1666464484
transform 1 0 14352 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_151
timestamp 1666464484
transform 1 0 14996 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_163
timestamp 1666464484
transform 1 0 16100 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_175
timestamp 1666464484
transform 1 0 17204 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_187
timestamp 1666464484
transform 1 0 18308 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_194
timestamp 1666464484
transform 1 0 18952 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_206
timestamp 1666464484
transform 1 0 20056 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_218
timestamp 1666464484
transform 1 0 21160 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_230
timestamp 1666464484
transform 1 0 22264 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_237
timestamp 1666464484
transform 1 0 22908 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_249
timestamp 1666464484
transform 1 0 24012 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_253
timestamp 1666464484
transform 1 0 24380 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_256
timestamp 1666464484
transform 1 0 24656 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_96_267
timestamp 1666464484
transform 1 0 25668 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_277
timestamp 1666464484
transform 1 0 26588 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_96_280
timestamp 1666464484
transform 1 0 26864 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_286
timestamp 1666464484
transform 1 0 27416 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_290
timestamp 1666464484
transform 1 0 27784 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_297
timestamp 1666464484
transform 1 0 28428 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_308
timestamp 1666464484
transform 1 0 29440 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_314
timestamp 1666464484
transform 1 0 29992 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_320
timestamp 1666464484
transform 1 0 30544 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_323
timestamp 1666464484
transform 1 0 30820 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_332
timestamp 1666464484
transform 1 0 31648 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_336
timestamp 1666464484
transform 1 0 32016 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_344
timestamp 1666464484
transform 1 0 32752 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_350
timestamp 1666464484
transform 1 0 33304 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_96_362
timestamp 1666464484
transform 1 0 34408 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_366
timestamp 1666464484
transform 1 0 34776 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_374
timestamp 1666464484
transform 1 0 35512 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_381
timestamp 1666464484
transform 1 0 36156 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_388
timestamp 1666464484
transform 1 0 36800 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_395
timestamp 1666464484
transform 1 0 37444 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_96_406
timestamp 1666464484
transform 1 0 38456 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_409
timestamp 1666464484
transform 1 0 38732 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_416
timestamp 1666464484
transform 1 0 39376 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_425
timestamp 1666464484
transform 1 0 40204 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_96_438
timestamp 1666464484
transform 1 0 41400 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_96_448
timestamp 1666464484
transform 1 0 42320 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_452
timestamp 1666464484
transform 1 0 42688 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_457
timestamp 1666464484
transform 1 0 43148 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_463
timestamp 1666464484
transform 1 0 43700 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_475
timestamp 1666464484
transform 1 0 44804 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_487
timestamp 1666464484
transform 1 0 45908 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_493
timestamp 1666464484
transform 1 0 46460 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_495
timestamp 1666464484
transform 1 0 46644 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_507
timestamp 1666464484
transform 1 0 47748 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_519
timestamp 1666464484
transform 1 0 48852 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_531
timestamp 1666464484
transform 1 0 49956 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_538
timestamp 1666464484
transform 1 0 50600 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_550
timestamp 1666464484
transform 1 0 51704 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_562
timestamp 1666464484
transform 1 0 52808 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_574
timestamp 1666464484
transform 1 0 53912 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_581
timestamp 1666464484
transform 1 0 54556 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_593
timestamp 1666464484
transform 1 0 55660 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_605
timestamp 1666464484
transform 1 0 56764 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_617
timestamp 1666464484
transform 1 0 57868 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_624
timestamp 1666464484
transform 1 0 58512 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1666464484
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1666464484
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1666464484
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_39
timestamp 1666464484
transform 1 0 4692 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_44
timestamp 1666464484
transform 1 0 5152 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_56
timestamp 1666464484
transform 1 0 6256 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_68
timestamp 1666464484
transform 1 0 7360 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_80
timestamp 1666464484
transform 1 0 8464 0 -1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_97_87
timestamp 1666464484
transform 1 0 9108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_99
timestamp 1666464484
transform 1 0 10212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_111
timestamp 1666464484
transform 1 0 11316 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_123
timestamp 1666464484
transform 1 0 12420 0 -1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_97_130
timestamp 1666464484
transform 1 0 13064 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_142
timestamp 1666464484
transform 1 0 14168 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_154
timestamp 1666464484
transform 1 0 15272 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_166
timestamp 1666464484
transform 1 0 16376 0 -1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_97_173
timestamp 1666464484
transform 1 0 17020 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_185
timestamp 1666464484
transform 1 0 18124 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_197
timestamp 1666464484
transform 1 0 19228 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_209
timestamp 1666464484
transform 1 0 20332 0 -1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_97_216
timestamp 1666464484
transform 1 0 20976 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_228
timestamp 1666464484
transform 1 0 22080 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_240
timestamp 1666464484
transform 1 0 23184 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_97_250
timestamp 1666464484
transform 1 0 24104 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_256
timestamp 1666464484
transform 1 0 24656 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_259
timestamp 1666464484
transform 1 0 24932 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_266
timestamp 1666464484
transform 1 0 25576 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_273
timestamp 1666464484
transform 1 0 26220 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_280
timestamp 1666464484
transform 1 0 26864 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_288
timestamp 1666464484
transform 1 0 27600 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_292
timestamp 1666464484
transform 1 0 27968 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_299
timestamp 1666464484
transform 1 0 28612 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_302
timestamp 1666464484
transform 1 0 28888 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_313
timestamp 1666464484
transform 1 0 29900 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_320
timestamp 1666464484
transform 1 0 30544 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1666464484
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_97_341
timestamp 1666464484
transform 1 0 32476 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_345
timestamp 1666464484
transform 1 0 32844 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_97_353
timestamp 1666464484
transform 1 0 33580 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_361
timestamp 1666464484
transform 1 0 34316 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_369
timestamp 1666464484
transform 1 0 35052 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_377
timestamp 1666464484
transform 1 0 35788 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_97_384
timestamp 1666464484
transform 1 0 36432 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_388
timestamp 1666464484
transform 1 0 36800 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_396
timestamp 1666464484
transform 1 0 37536 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_406
timestamp 1666464484
transform 1 0 38456 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_417
timestamp 1666464484
transform 1 0 39468 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_421
timestamp 1666464484
transform 1 0 39836 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_428
timestamp 1666464484
transform 1 0 40480 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_431
timestamp 1666464484
transform 1 0 40756 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_438
timestamp 1666464484
transform 1 0 41400 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_450
timestamp 1666464484
transform 1 0 42504 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_461
timestamp 1666464484
transform 1 0 43516 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_471
timestamp 1666464484
transform 1 0 44436 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_474
timestamp 1666464484
transform 1 0 44712 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_479
timestamp 1666464484
transform 1 0 45172 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_485
timestamp 1666464484
transform 1 0 45724 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_491
timestamp 1666464484
transform 1 0 46276 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_503
timestamp 1666464484
transform 1 0 47380 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_515
timestamp 1666464484
transform 1 0 48484 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1666464484
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1666464484
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1666464484
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1666464484
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_97_560
timestamp 1666464484
transform 1 0 52624 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_572
timestamp 1666464484
transform 1 0 53728 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_584
timestamp 1666464484
transform 1 0 54832 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_596
timestamp 1666464484
transform 1 0 55936 0 -1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_97_603
timestamp 1666464484
transform 1 0 56580 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_615
timestamp 1666464484
transform 1 0 57684 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_623
timestamp 1666464484
transform 1 0 58420 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1666464484
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_15
timestamp 1666464484
transform 1 0 2484 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_22
timestamp 1666464484
transform 1 0 3128 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_34
timestamp 1666464484
transform 1 0 4232 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_46
timestamp 1666464484
transform 1 0 5336 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_58
timestamp 1666464484
transform 1 0 6440 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1666464484
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_77
timestamp 1666464484
transform 1 0 8188 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_89
timestamp 1666464484
transform 1 0 9292 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_101
timestamp 1666464484
transform 1 0 10396 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_108
timestamp 1666464484
transform 1 0 11040 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_120
timestamp 1666464484
transform 1 0 12144 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_132
timestamp 1666464484
transform 1 0 13248 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_144
timestamp 1666464484
transform 1 0 14352 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_151
timestamp 1666464484
transform 1 0 14996 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_163
timestamp 1666464484
transform 1 0 16100 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_175
timestamp 1666464484
transform 1 0 17204 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_187
timestamp 1666464484
transform 1 0 18308 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_194
timestamp 1666464484
transform 1 0 18952 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_206
timestamp 1666464484
transform 1 0 20056 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_218
timestamp 1666464484
transform 1 0 21160 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_230
timestamp 1666464484
transform 1 0 22264 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_98_237
timestamp 1666464484
transform 1 0 22908 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_241
timestamp 1666464484
transform 1 0 23276 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_244
timestamp 1666464484
transform 1 0 23552 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_251
timestamp 1666464484
transform 1 0 24196 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_258
timestamp 1666464484
transform 1 0 24840 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_265
timestamp 1666464484
transform 1 0 25484 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_273
timestamp 1666464484
transform 1 0 26220 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_98_280
timestamp 1666464484
transform 1 0 26864 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_286
timestamp 1666464484
transform 1 0 27416 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_295
timestamp 1666464484
transform 1 0 28244 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_306
timestamp 1666464484
transform 1 0 29256 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_314
timestamp 1666464484
transform 1 0 29992 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_320
timestamp 1666464484
transform 1 0 30544 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_323
timestamp 1666464484
transform 1 0 30820 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_333
timestamp 1666464484
transform 1 0 31740 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_343
timestamp 1666464484
transform 1 0 32660 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_353
timestamp 1666464484
transform 1 0 33580 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_357
timestamp 1666464484
transform 1 0 33948 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_363
timestamp 1666464484
transform 1 0 34500 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_366
timestamp 1666464484
transform 1 0 34776 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_98_375
timestamp 1666464484
transform 1 0 35604 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_98_389
timestamp 1666464484
transform 1 0 36892 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_395
timestamp 1666464484
transform 1 0 37444 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_406
timestamp 1666464484
transform 1 0 38456 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_409
timestamp 1666464484
transform 1 0 38732 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_416
timestamp 1666464484
transform 1 0 39376 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_423
timestamp 1666464484
transform 1 0 40020 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_433
timestamp 1666464484
transform 1 0 40940 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_443
timestamp 1666464484
transform 1 0 41860 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_449
timestamp 1666464484
transform 1 0 42412 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_98_452
timestamp 1666464484
transform 1 0 42688 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_98_465
timestamp 1666464484
transform 1 0 43884 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_473
timestamp 1666464484
transform 1 0 44620 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_480
timestamp 1666464484
transform 1 0 45264 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_487
timestamp 1666464484
transform 1 0 45908 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_493
timestamp 1666464484
transform 1 0 46460 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_495
timestamp 1666464484
transform 1 0 46644 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_98_499
timestamp 1666464484
transform 1 0 47012 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_98_507
timestamp 1666464484
transform 1 0 47748 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_511
timestamp 1666464484
transform 1 0 48116 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_514
timestamp 1666464484
transform 1 0 48392 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_526
timestamp 1666464484
transform 1 0 49496 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_534
timestamp 1666464484
transform 1 0 50232 0 1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_98_538
timestamp 1666464484
transform 1 0 50600 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_550
timestamp 1666464484
transform 1 0 51704 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_562
timestamp 1666464484
transform 1 0 52808 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_574
timestamp 1666464484
transform 1 0 53912 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_581
timestamp 1666464484
transform 1 0 54556 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_593
timestamp 1666464484
transform 1 0 55660 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_605
timestamp 1666464484
transform 1 0 56764 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_617
timestamp 1666464484
transform 1 0 57868 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_624
timestamp 1666464484
transform 1 0 58512 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1666464484
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1666464484
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1666464484
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_39
timestamp 1666464484
transform 1 0 4692 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_44
timestamp 1666464484
transform 1 0 5152 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_56
timestamp 1666464484
transform 1 0 6256 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_68
timestamp 1666464484
transform 1 0 7360 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_80
timestamp 1666464484
transform 1 0 8464 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_87
timestamp 1666464484
transform 1 0 9108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_99
timestamp 1666464484
transform 1 0 10212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_111
timestamp 1666464484
transform 1 0 11316 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_123
timestamp 1666464484
transform 1 0 12420 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_130
timestamp 1666464484
transform 1 0 13064 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_142
timestamp 1666464484
transform 1 0 14168 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_154
timestamp 1666464484
transform 1 0 15272 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_166
timestamp 1666464484
transform 1 0 16376 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_173
timestamp 1666464484
transform 1 0 17020 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_185
timestamp 1666464484
transform 1 0 18124 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_197
timestamp 1666464484
transform 1 0 19228 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_209
timestamp 1666464484
transform 1 0 20332 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_216
timestamp 1666464484
transform 1 0 20976 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_228
timestamp 1666464484
transform 1 0 22080 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_99_237
timestamp 1666464484
transform 1 0 22908 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_241
timestamp 1666464484
transform 1 0 23276 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_245
timestamp 1666464484
transform 1 0 23644 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_254
timestamp 1666464484
transform 1 0 24472 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_99_259
timestamp 1666464484
transform 1 0 24932 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_267
timestamp 1666464484
transform 1 0 25668 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_277
timestamp 1666464484
transform 1 0 26588 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_286
timestamp 1666464484
transform 1 0 27416 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_292
timestamp 1666464484
transform 1 0 27968 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_99_298
timestamp 1666464484
transform 1 0 28520 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_99_302
timestamp 1666464484
transform 1 0 28888 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_99_313
timestamp 1666464484
transform 1 0 29900 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_321
timestamp 1666464484
transform 1 0 30636 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1666464484
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1666464484
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_342
timestamp 1666464484
transform 1 0 32568 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_345
timestamp 1666464484
transform 1 0 32844 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_353
timestamp 1666464484
transform 1 0 33580 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_363
timestamp 1666464484
transform 1 0 34500 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_369
timestamp 1666464484
transform 1 0 35052 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_381
timestamp 1666464484
transform 1 0 36156 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_99_388
timestamp 1666464484
transform 1 0 36800 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_397
timestamp 1666464484
transform 1 0 37628 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_407
timestamp 1666464484
transform 1 0 38548 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_414
timestamp 1666464484
transform 1 0 39192 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_426
timestamp 1666464484
transform 1 0 40296 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_431
timestamp 1666464484
transform 1 0 40756 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_439
timestamp 1666464484
transform 1 0 41492 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_449
timestamp 1666464484
transform 1 0 42412 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_453
timestamp 1666464484
transform 1 0 42780 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_461
timestamp 1666464484
transform 1 0 43516 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_471
timestamp 1666464484
transform 1 0 44436 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_474
timestamp 1666464484
transform 1 0 44712 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_481
timestamp 1666464484
transform 1 0 45356 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_488
timestamp 1666464484
transform 1 0 46000 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_495
timestamp 1666464484
transform 1 0 46644 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_502
timestamp 1666464484
transform 1 0 47288 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_509
timestamp 1666464484
transform 1 0 47932 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_515
timestamp 1666464484
transform 1 0 48484 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_517
timestamp 1666464484
transform 1 0 48668 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_522
timestamp 1666464484
transform 1 0 49128 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_529
timestamp 1666464484
transform 1 0 49772 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_535
timestamp 1666464484
transform 1 0 50324 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_549
timestamp 1666464484
transform 1 0 51612 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_557
timestamp 1666464484
transform 1 0 52348 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_560
timestamp 1666464484
transform 1 0 52624 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_99_564
timestamp 1666464484
transform 1 0 52992 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_574
timestamp 1666464484
transform 1 0 53912 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_586
timestamp 1666464484
transform 1 0 55016 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_598
timestamp 1666464484
transform 1 0 56120 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_603
timestamp 1666464484
transform 1 0 56580 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_615
timestamp 1666464484
transform 1 0 57684 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_623
timestamp 1666464484
transform 1 0 58420 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1666464484
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_15
timestamp 1666464484
transform 1 0 2484 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_100_22
timestamp 1666464484
transform 1 0 3128 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_26
timestamp 1666464484
transform 1 0 3496 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1666464484
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1666464484
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_53
timestamp 1666464484
transform 1 0 5980 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_57
timestamp 1666464484
transform 1 0 6348 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_63
timestamp 1666464484
transform 1 0 6900 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_65
timestamp 1666464484
transform 1 0 7084 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_72
timestamp 1666464484
transform 1 0 7728 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_84
timestamp 1666464484
transform 1 0 8832 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_96
timestamp 1666464484
transform 1 0 9936 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_104
timestamp 1666464484
transform 1 0 10672 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_100_108
timestamp 1666464484
transform 1 0 11040 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_100_117
timestamp 1666464484
transform 1 0 11868 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_123
timestamp 1666464484
transform 1 0 12420 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_132
timestamp 1666464484
transform 1 0 13248 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_144
timestamp 1666464484
transform 1 0 14352 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_151
timestamp 1666464484
transform 1 0 14996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_163
timestamp 1666464484
transform 1 0 16100 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_171
timestamp 1666464484
transform 1 0 16836 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1666464484
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_189
timestamp 1666464484
transform 1 0 18492 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_194
timestamp 1666464484
transform 1 0 18952 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_199
timestamp 1666464484
transform 1 0 19412 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_211
timestamp 1666464484
transform 1 0 20516 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_100_222
timestamp 1666464484
transform 1 0 21528 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_230
timestamp 1666464484
transform 1 0 22264 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_234
timestamp 1666464484
transform 1 0 22632 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_237
timestamp 1666464484
transform 1 0 22908 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_241
timestamp 1666464484
transform 1 0 23276 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_253
timestamp 1666464484
transform 1 0 24380 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_259
timestamp 1666464484
transform 1 0 24932 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_268
timestamp 1666464484
transform 1 0 25760 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_277
timestamp 1666464484
transform 1 0 26588 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_280
timestamp 1666464484
transform 1 0 26864 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_290
timestamp 1666464484
transform 1 0 27784 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_301
timestamp 1666464484
transform 1 0 28796 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_314
timestamp 1666464484
transform 1 0 29992 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_320
timestamp 1666464484
transform 1 0 30544 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_323
timestamp 1666464484
transform 1 0 30820 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_328
timestamp 1666464484
transform 1 0 31280 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_340
timestamp 1666464484
transform 1 0 32384 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_348
timestamp 1666464484
transform 1 0 33120 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_356
timestamp 1666464484
transform 1 0 33856 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_363
timestamp 1666464484
transform 1 0 34500 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_366
timestamp 1666464484
transform 1 0 34776 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_375
timestamp 1666464484
transform 1 0 35604 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_389
timestamp 1666464484
transform 1 0 36892 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_395
timestamp 1666464484
transform 1 0 37444 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_406
timestamp 1666464484
transform 1 0 38456 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_409
timestamp 1666464484
transform 1 0 38732 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_100_421
timestamp 1666464484
transform 1 0 39836 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_427
timestamp 1666464484
transform 1 0 40388 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_436
timestamp 1666464484
transform 1 0 41216 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_447
timestamp 1666464484
transform 1 0 42228 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_452
timestamp 1666464484
transform 1 0 42688 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_460
timestamp 1666464484
transform 1 0 43424 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_464
timestamp 1666464484
transform 1 0 43792 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_475
timestamp 1666464484
transform 1 0 44804 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_482
timestamp 1666464484
transform 1 0 45448 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_489
timestamp 1666464484
transform 1 0 46092 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_493
timestamp 1666464484
transform 1 0 46460 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_495
timestamp 1666464484
transform 1 0 46644 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_500
timestamp 1666464484
transform 1 0 47104 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_507
timestamp 1666464484
transform 1 0 47748 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_513
timestamp 1666464484
transform 1 0 48300 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_524
timestamp 1666464484
transform 1 0 49312 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_531
timestamp 1666464484
transform 1 0 49956 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_100_538
timestamp 1666464484
transform 1 0 50600 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_543
timestamp 1666464484
transform 1 0 51060 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_550
timestamp 1666464484
transform 1 0 51704 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_557
timestamp 1666464484
transform 1 0 52348 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_564
timestamp 1666464484
transform 1 0 52992 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_571
timestamp 1666464484
transform 1 0 53636 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_578
timestamp 1666464484
transform 1 0 54280 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_100_581
timestamp 1666464484
transform 1 0 54556 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_587
timestamp 1666464484
transform 1 0 55108 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_593
timestamp 1666464484
transform 1 0 55660 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_602
timestamp 1666464484
transform 1 0 56488 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_614
timestamp 1666464484
transform 1 0 57592 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_622
timestamp 1666464484
transform 1 0 58328 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_100_624
timestamp 1666464484
transform 1 0 58512 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1666464484
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_15
timestamp 1666464484
transform 1 0 2484 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_101_22
timestamp 1666464484
transform 1 0 3128 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_28
timestamp 1666464484
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_33
timestamp 1666464484
transform 1 0 4140 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_40
timestamp 1666464484
transform 1 0 4784 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_43
timestamp 1666464484
transform 1 0 5060 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_49
timestamp 1666464484
transform 1 0 5612 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_57
timestamp 1666464484
transform 1 0 6348 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_61
timestamp 1666464484
transform 1 0 6716 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_64
timestamp 1666464484
transform 1 0 6992 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_68
timestamp 1666464484
transform 1 0 7360 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_75
timestamp 1666464484
transform 1 0 8004 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_82
timestamp 1666464484
transform 1 0 8648 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_85
timestamp 1666464484
transform 1 0 8924 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_92
timestamp 1666464484
transform 1 0 9568 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_98
timestamp 1666464484
transform 1 0 10120 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_102
timestamp 1666464484
transform 1 0 10488 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_106
timestamp 1666464484
transform 1 0 10856 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_112
timestamp 1666464484
transform 1 0 11408 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_118
timestamp 1666464484
transform 1 0 11960 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_123
timestamp 1666464484
transform 1 0 12420 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_127
timestamp 1666464484
transform 1 0 12788 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_133
timestamp 1666464484
transform 1 0 13340 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_138
timestamp 1666464484
transform 1 0 13800 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_145
timestamp 1666464484
transform 1 0 14444 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_148
timestamp 1666464484
transform 1 0 14720 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_154
timestamp 1666464484
transform 1 0 15272 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_158
timestamp 1666464484
transform 1 0 15640 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_162
timestamp 1666464484
transform 1 0 16008 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_101_169
timestamp 1666464484
transform 1 0 16652 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_175
timestamp 1666464484
transform 1 0 17204 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_183
timestamp 1666464484
transform 1 0 17940 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_190
timestamp 1666464484
transform 1 0 18584 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_198
timestamp 1666464484
transform 1 0 19320 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_101_207
timestamp 1666464484
transform 1 0 20148 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_211
timestamp 1666464484
transform 1 0 20516 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_217
timestamp 1666464484
transform 1 0 21068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_223
timestamp 1666464484
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_228
timestamp 1666464484
transform 1 0 22080 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_232
timestamp 1666464484
transform 1 0 22448 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_242
timestamp 1666464484
transform 1 0 23368 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_250
timestamp 1666464484
transform 1 0 24104 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_253
timestamp 1666464484
transform 1 0 24380 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_260
timestamp 1666464484
transform 1 0 25024 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_269
timestamp 1666464484
transform 1 0 25852 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_274
timestamp 1666464484
transform 1 0 26312 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_284
timestamp 1666464484
transform 1 0 27232 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_292
timestamp 1666464484
transform 1 0 27968 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_295
timestamp 1666464484
transform 1 0 28244 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_301
timestamp 1666464484
transform 1 0 28796 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_310
timestamp 1666464484
transform 1 0 29624 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_314
timestamp 1666464484
transform 1 0 29992 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_316
timestamp 1666464484
transform 1 0 30176 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_322
timestamp 1666464484
transform 1 0 30728 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_326
timestamp 1666464484
transform 1 0 31096 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_333
timestamp 1666464484
transform 1 0 31740 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_337
timestamp 1666464484
transform 1 0 32108 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_349
timestamp 1666464484
transform 1 0 33212 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_355
timestamp 1666464484
transform 1 0 33764 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_358
timestamp 1666464484
transform 1 0 34040 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_368
timestamp 1666464484
transform 1 0 34960 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_101_375
timestamp 1666464484
transform 1 0 35604 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_379
timestamp 1666464484
transform 1 0 35972 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_391
timestamp 1666464484
transform 1 0 37076 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_397
timestamp 1666464484
transform 1 0 37628 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_400
timestamp 1666464484
transform 1 0 37904 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_412
timestamp 1666464484
transform 1 0 39008 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_418
timestamp 1666464484
transform 1 0 39560 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_421
timestamp 1666464484
transform 1 0 39836 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_430
timestamp 1666464484
transform 1 0 40664 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_439
timestamp 1666464484
transform 1 0 41492 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_442
timestamp 1666464484
transform 1 0 41768 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_446
timestamp 1666464484
transform 1 0 42136 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_460
timestamp 1666464484
transform 1 0 43424 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_463
timestamp 1666464484
transform 1 0 43700 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_471
timestamp 1666464484
transform 1 0 44436 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_478
timestamp 1666464484
transform 1 0 45080 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_482
timestamp 1666464484
transform 1 0 45448 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_484
timestamp 1666464484
transform 1 0 45632 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_490
timestamp 1666464484
transform 1 0 46184 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_497
timestamp 1666464484
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1666464484
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_505
timestamp 1666464484
transform 1 0 47564 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_517
timestamp 1666464484
transform 1 0 48668 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_523
timestamp 1666464484
transform 1 0 49220 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_101_526
timestamp 1666464484
transform 1 0 49496 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_539
timestamp 1666464484
transform 1 0 50692 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_545
timestamp 1666464484
transform 1 0 51244 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_547
timestamp 1666464484
transform 1 0 51428 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_553
timestamp 1666464484
transform 1 0 51980 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_101_565
timestamp 1666464484
transform 1 0 53084 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_568
timestamp 1666464484
transform 1 0 53360 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_578
timestamp 1666464484
transform 1 0 54280 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_101_585
timestamp 1666464484
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_589
timestamp 1666464484
transform 1 0 55292 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_595
timestamp 1666464484
transform 1 0 55844 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_602
timestamp 1666464484
transform 1 0 56488 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_608
timestamp 1666464484
transform 1 0 57040 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_610
timestamp 1666464484
transform 1 0 57224 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_622
timestamp 1666464484
transform 1 0 58328 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666464484
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666464484
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666464484
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666464484
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666464484
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666464484
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666464484
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666464484
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666464484
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666464484
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666464484
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666464484
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666464484
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666464484
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666464484
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666464484
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666464484
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666464484
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666464484
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666464484
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666464484
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666464484
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666464484
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666464484
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666464484
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666464484
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666464484
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666464484
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666464484
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666464484
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666464484
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666464484
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666464484
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666464484
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666464484
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666464484
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1666464484
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1666464484
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1666464484
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1666464484
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1666464484
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1666464484
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1666464484
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1666464484
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1666464484
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1666464484
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1666464484
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1666464484
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1666464484
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1666464484
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1666464484
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1666464484
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1666464484
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1666464484
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1666464484
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1666464484
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1666464484
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1666464484
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1666464484
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1666464484
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1666464484
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1666464484
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1666464484
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1666464484
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1666464484
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1666464484
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1666464484
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1666464484
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1666464484
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1666464484
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1666464484
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1666464484
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1666464484
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1666464484
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 4968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 10764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 12696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 14628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 20424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 22356 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 26220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 28152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 30084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 33948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 35880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 37812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 41676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 43608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 45540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 49404 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 51336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 53268 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 57132 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 5060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 9016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 12972 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 16928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 20884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 24840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 28796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 32752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 36708 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 40664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 44620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 48576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 56488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 3036 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 6992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 10948 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 14904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 18860 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 22816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 26772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 30728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 34684 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 38640 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 42596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 46552 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 50508 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 54464 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 58420 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 5060 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 9016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 12972 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 16928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 20884 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 24840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 28796 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 32752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 36708 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 40664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 44620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 48576 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 56488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 3036 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 6992 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 10948 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 14904 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 18860 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 22816 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 26772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 30728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 34684 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 38640 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 42596 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 46552 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 50508 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 54464 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 58420 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 9016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 12972 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 16928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 20884 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 24840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 28796 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 32752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 36708 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 40664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 44620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 48576 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 56488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 6992 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 10948 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 14904 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 18860 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 22816 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 26772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 30728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 34684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 38640 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 42596 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 46552 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 50508 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 54464 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 58420 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 5060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 9016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 12972 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 16928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 20884 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 24840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 28796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 32752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 36708 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 40664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 44620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 48576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 56488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 3036 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 6992 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 10948 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 14904 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 18860 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 22816 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 26772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 30728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 34684 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 38640 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 42596 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 46552 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 50508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 54464 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 58420 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 5060 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 9016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 12972 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 16928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 20884 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 24840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 28796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 32752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 36708 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 40664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 44620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 48576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 56488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 3036 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 6992 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 10948 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 14904 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 18860 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 22816 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 26772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 30728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 34684 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 38640 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 42596 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 46552 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 50508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 54464 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 58420 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 5060 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 9016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 12972 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 16928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 20884 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 24840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 28796 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 32752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 36708 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 40664 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 44620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 48576 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 56488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 3036 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 6992 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 10948 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 14904 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 18860 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 22816 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 26772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 30728 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 34684 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 38640 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 42596 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 46552 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 50508 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 54464 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 58420 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 5060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 9016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 12972 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 16928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 20884 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 24840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 28796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 32752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 36708 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 40664 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 44620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 48576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 56488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 3036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 6992 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 10948 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 14904 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 18860 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 22816 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 26772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 30728 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 34684 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 38640 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 42596 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 46552 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 50508 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 54464 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 58420 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 5060 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 9016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 12972 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 16928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 20884 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 24840 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 28796 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 32752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 36708 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 40664 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 44620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 48576 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 56488 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 3036 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 6992 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 10948 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 14904 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 18860 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 22816 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 26772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 30728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 34684 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 38640 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 42596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 46552 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 50508 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 54464 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 58420 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 9016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 12972 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 16928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 20884 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 24840 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 28796 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 32752 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 36708 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 40664 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 44620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 48576 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 56488 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 3036 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 6992 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 10948 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 14904 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 18860 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 22816 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 26772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 30728 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 34684 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 38640 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 42596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 46552 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 50508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 54464 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 58420 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 5060 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 9016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 16928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 20884 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 24840 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 28796 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 32752 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 36708 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 40664 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 44620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 48576 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 56488 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 3036 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 6992 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 10948 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 14904 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 18860 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 22816 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 26772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 30728 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 34684 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 38640 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 42596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 46552 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 50508 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 54464 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 58420 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 5060 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 9016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 12972 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 16928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 20884 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 24840 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 28796 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 32752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 36708 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 40664 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 44620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 48576 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 56488 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 3036 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 6992 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 10948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 14904 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 18860 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 22816 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 26772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 30728 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 34684 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 38640 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 42596 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 46552 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 50508 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 54464 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 58420 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 5060 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 9016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 12972 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 16928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 20884 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 24840 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 28796 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 32752 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 36708 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 40664 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 44620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 48576 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666464484
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666464484
transform 1 0 56488 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666464484
transform 1 0 3036 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666464484
transform 1 0 6992 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666464484
transform 1 0 10948 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666464484
transform 1 0 14904 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666464484
transform 1 0 18860 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666464484
transform 1 0 22816 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666464484
transform 1 0 26772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666464484
transform 1 0 30728 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666464484
transform 1 0 34684 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666464484
transform 1 0 38640 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666464484
transform 1 0 42596 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666464484
transform 1 0 46552 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666464484
transform 1 0 50508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666464484
transform 1 0 54464 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666464484
transform 1 0 58420 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666464484
transform 1 0 5060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666464484
transform 1 0 9016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666464484
transform 1 0 12972 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666464484
transform 1 0 16928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666464484
transform 1 0 20884 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666464484
transform 1 0 24840 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666464484
transform 1 0 28796 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666464484
transform 1 0 32752 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666464484
transform 1 0 36708 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666464484
transform 1 0 40664 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666464484
transform 1 0 44620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666464484
transform 1 0 48576 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666464484
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666464484
transform 1 0 56488 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666464484
transform 1 0 3036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666464484
transform 1 0 6992 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666464484
transform 1 0 10948 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666464484
transform 1 0 14904 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666464484
transform 1 0 18860 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666464484
transform 1 0 22816 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666464484
transform 1 0 26772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666464484
transform 1 0 30728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666464484
transform 1 0 34684 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666464484
transform 1 0 38640 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666464484
transform 1 0 42596 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666464484
transform 1 0 46552 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666464484
transform 1 0 50508 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666464484
transform 1 0 54464 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666464484
transform 1 0 58420 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666464484
transform 1 0 5060 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666464484
transform 1 0 9016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666464484
transform 1 0 12972 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666464484
transform 1 0 16928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666464484
transform 1 0 20884 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666464484
transform 1 0 24840 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666464484
transform 1 0 28796 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666464484
transform 1 0 32752 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666464484
transform 1 0 36708 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666464484
transform 1 0 40664 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666464484
transform 1 0 44620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666464484
transform 1 0 48576 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666464484
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666464484
transform 1 0 56488 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666464484
transform 1 0 3036 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666464484
transform 1 0 6992 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666464484
transform 1 0 10948 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666464484
transform 1 0 14904 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666464484
transform 1 0 18860 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666464484
transform 1 0 22816 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666464484
transform 1 0 26772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666464484
transform 1 0 30728 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666464484
transform 1 0 34684 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666464484
transform 1 0 38640 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666464484
transform 1 0 42596 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666464484
transform 1 0 46552 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666464484
transform 1 0 50508 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666464484
transform 1 0 54464 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666464484
transform 1 0 58420 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666464484
transform 1 0 5060 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666464484
transform 1 0 9016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666464484
transform 1 0 12972 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666464484
transform 1 0 16928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666464484
transform 1 0 20884 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666464484
transform 1 0 24840 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666464484
transform 1 0 28796 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666464484
transform 1 0 32752 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666464484
transform 1 0 36708 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666464484
transform 1 0 40664 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666464484
transform 1 0 44620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666464484
transform 1 0 48576 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666464484
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666464484
transform 1 0 56488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666464484
transform 1 0 3036 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666464484
transform 1 0 6992 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666464484
transform 1 0 10948 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666464484
transform 1 0 14904 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666464484
transform 1 0 18860 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666464484
transform 1 0 22816 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666464484
transform 1 0 26772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666464484
transform 1 0 30728 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666464484
transform 1 0 34684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666464484
transform 1 0 38640 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666464484
transform 1 0 42596 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666464484
transform 1 0 46552 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666464484
transform 1 0 50508 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666464484
transform 1 0 54464 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666464484
transform 1 0 58420 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666464484
transform 1 0 5060 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666464484
transform 1 0 9016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666464484
transform 1 0 12972 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666464484
transform 1 0 16928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666464484
transform 1 0 20884 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666464484
transform 1 0 24840 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666464484
transform 1 0 28796 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666464484
transform 1 0 32752 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666464484
transform 1 0 36708 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666464484
transform 1 0 40664 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666464484
transform 1 0 44620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666464484
transform 1 0 48576 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666464484
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666464484
transform 1 0 56488 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666464484
transform 1 0 3036 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666464484
transform 1 0 6992 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666464484
transform 1 0 10948 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666464484
transform 1 0 14904 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666464484
transform 1 0 18860 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666464484
transform 1 0 22816 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666464484
transform 1 0 26772 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666464484
transform 1 0 30728 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666464484
transform 1 0 34684 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666464484
transform 1 0 38640 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666464484
transform 1 0 42596 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666464484
transform 1 0 46552 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666464484
transform 1 0 50508 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666464484
transform 1 0 54464 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666464484
transform 1 0 58420 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666464484
transform 1 0 5060 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666464484
transform 1 0 9016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666464484
transform 1 0 12972 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666464484
transform 1 0 16928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666464484
transform 1 0 20884 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666464484
transform 1 0 24840 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666464484
transform 1 0 28796 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666464484
transform 1 0 32752 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666464484
transform 1 0 36708 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666464484
transform 1 0 40664 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666464484
transform 1 0 44620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666464484
transform 1 0 48576 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666464484
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666464484
transform 1 0 56488 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666464484
transform 1 0 3036 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666464484
transform 1 0 6992 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666464484
transform 1 0 10948 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666464484
transform 1 0 14904 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666464484
transform 1 0 18860 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666464484
transform 1 0 22816 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666464484
transform 1 0 26772 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666464484
transform 1 0 30728 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666464484
transform 1 0 34684 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666464484
transform 1 0 38640 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666464484
transform 1 0 42596 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666464484
transform 1 0 46552 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666464484
transform 1 0 50508 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666464484
transform 1 0 54464 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666464484
transform 1 0 58420 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666464484
transform 1 0 5060 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666464484
transform 1 0 9016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666464484
transform 1 0 12972 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666464484
transform 1 0 16928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666464484
transform 1 0 20884 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666464484
transform 1 0 24840 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666464484
transform 1 0 28796 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666464484
transform 1 0 32752 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666464484
transform 1 0 36708 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666464484
transform 1 0 40664 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666464484
transform 1 0 44620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666464484
transform 1 0 48576 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666464484
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666464484
transform 1 0 56488 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666464484
transform 1 0 3036 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666464484
transform 1 0 6992 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666464484
transform 1 0 10948 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666464484
transform 1 0 14904 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666464484
transform 1 0 18860 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666464484
transform 1 0 22816 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666464484
transform 1 0 26772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666464484
transform 1 0 30728 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666464484
transform 1 0 34684 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666464484
transform 1 0 38640 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666464484
transform 1 0 42596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666464484
transform 1 0 46552 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666464484
transform 1 0 50508 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666464484
transform 1 0 54464 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666464484
transform 1 0 58420 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666464484
transform 1 0 5060 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666464484
transform 1 0 9016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666464484
transform 1 0 12972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666464484
transform 1 0 16928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666464484
transform 1 0 20884 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666464484
transform 1 0 24840 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666464484
transform 1 0 28796 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666464484
transform 1 0 32752 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666464484
transform 1 0 36708 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666464484
transform 1 0 40664 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666464484
transform 1 0 44620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666464484
transform 1 0 48576 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666464484
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666464484
transform 1 0 56488 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666464484
transform 1 0 3036 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666464484
transform 1 0 6992 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666464484
transform 1 0 10948 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666464484
transform 1 0 14904 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666464484
transform 1 0 18860 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666464484
transform 1 0 22816 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666464484
transform 1 0 26772 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666464484
transform 1 0 30728 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666464484
transform 1 0 34684 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666464484
transform 1 0 38640 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666464484
transform 1 0 42596 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666464484
transform 1 0 46552 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666464484
transform 1 0 50508 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666464484
transform 1 0 54464 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666464484
transform 1 0 58420 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666464484
transform 1 0 5060 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666464484
transform 1 0 9016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666464484
transform 1 0 12972 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666464484
transform 1 0 16928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666464484
transform 1 0 20884 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666464484
transform 1 0 24840 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666464484
transform 1 0 28796 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666464484
transform 1 0 32752 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666464484
transform 1 0 36708 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666464484
transform 1 0 40664 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666464484
transform 1 0 44620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666464484
transform 1 0 48576 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666464484
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666464484
transform 1 0 56488 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666464484
transform 1 0 3036 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666464484
transform 1 0 6992 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666464484
transform 1 0 10948 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666464484
transform 1 0 14904 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666464484
transform 1 0 18860 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666464484
transform 1 0 22816 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666464484
transform 1 0 26772 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666464484
transform 1 0 30728 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666464484
transform 1 0 34684 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666464484
transform 1 0 38640 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666464484
transform 1 0 42596 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666464484
transform 1 0 46552 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666464484
transform 1 0 50508 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666464484
transform 1 0 54464 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666464484
transform 1 0 58420 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666464484
transform 1 0 5060 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666464484
transform 1 0 9016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666464484
transform 1 0 12972 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666464484
transform 1 0 16928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666464484
transform 1 0 20884 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666464484
transform 1 0 24840 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666464484
transform 1 0 28796 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666464484
transform 1 0 32752 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666464484
transform 1 0 36708 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666464484
transform 1 0 40664 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666464484
transform 1 0 44620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666464484
transform 1 0 48576 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666464484
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666464484
transform 1 0 56488 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666464484
transform 1 0 3036 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666464484
transform 1 0 6992 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666464484
transform 1 0 10948 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666464484
transform 1 0 14904 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666464484
transform 1 0 18860 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666464484
transform 1 0 22816 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666464484
transform 1 0 26772 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666464484
transform 1 0 30728 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666464484
transform 1 0 34684 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666464484
transform 1 0 38640 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666464484
transform 1 0 42596 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666464484
transform 1 0 46552 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666464484
transform 1 0 50508 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666464484
transform 1 0 54464 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666464484
transform 1 0 58420 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666464484
transform 1 0 5060 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666464484
transform 1 0 9016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666464484
transform 1 0 12972 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666464484
transform 1 0 16928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666464484
transform 1 0 20884 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666464484
transform 1 0 24840 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666464484
transform 1 0 28796 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666464484
transform 1 0 32752 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666464484
transform 1 0 36708 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666464484
transform 1 0 40664 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666464484
transform 1 0 44620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666464484
transform 1 0 48576 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666464484
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666464484
transform 1 0 56488 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666464484
transform 1 0 3036 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666464484
transform 1 0 6992 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666464484
transform 1 0 10948 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666464484
transform 1 0 14904 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666464484
transform 1 0 18860 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666464484
transform 1 0 22816 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666464484
transform 1 0 26772 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666464484
transform 1 0 30728 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666464484
transform 1 0 34684 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666464484
transform 1 0 38640 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666464484
transform 1 0 42596 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666464484
transform 1 0 46552 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666464484
transform 1 0 50508 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666464484
transform 1 0 54464 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666464484
transform 1 0 58420 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666464484
transform 1 0 5060 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666464484
transform 1 0 9016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666464484
transform 1 0 12972 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666464484
transform 1 0 16928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666464484
transform 1 0 20884 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666464484
transform 1 0 24840 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666464484
transform 1 0 28796 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666464484
transform 1 0 32752 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666464484
transform 1 0 36708 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666464484
transform 1 0 40664 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666464484
transform 1 0 44620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666464484
transform 1 0 48576 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666464484
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666464484
transform 1 0 56488 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666464484
transform 1 0 3036 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666464484
transform 1 0 6992 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666464484
transform 1 0 10948 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666464484
transform 1 0 14904 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666464484
transform 1 0 18860 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666464484
transform 1 0 22816 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666464484
transform 1 0 26772 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666464484
transform 1 0 30728 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666464484
transform 1 0 34684 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666464484
transform 1 0 38640 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666464484
transform 1 0 42596 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666464484
transform 1 0 46552 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666464484
transform 1 0 50508 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666464484
transform 1 0 54464 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666464484
transform 1 0 58420 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666464484
transform 1 0 5060 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666464484
transform 1 0 9016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666464484
transform 1 0 12972 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666464484
transform 1 0 16928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666464484
transform 1 0 20884 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666464484
transform 1 0 24840 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666464484
transform 1 0 28796 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666464484
transform 1 0 32752 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666464484
transform 1 0 36708 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666464484
transform 1 0 40664 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666464484
transform 1 0 44620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666464484
transform 1 0 48576 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666464484
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666464484
transform 1 0 56488 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666464484
transform 1 0 3036 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666464484
transform 1 0 6992 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666464484
transform 1 0 10948 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666464484
transform 1 0 14904 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666464484
transform 1 0 18860 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666464484
transform 1 0 22816 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666464484
transform 1 0 26772 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666464484
transform 1 0 30728 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666464484
transform 1 0 34684 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666464484
transform 1 0 38640 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666464484
transform 1 0 42596 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666464484
transform 1 0 46552 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666464484
transform 1 0 50508 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666464484
transform 1 0 54464 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666464484
transform 1 0 58420 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666464484
transform 1 0 5060 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666464484
transform 1 0 9016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1666464484
transform 1 0 12972 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1666464484
transform 1 0 16928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1666464484
transform 1 0 20884 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1666464484
transform 1 0 24840 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1666464484
transform 1 0 28796 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1666464484
transform 1 0 32752 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1666464484
transform 1 0 36708 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1666464484
transform 1 0 40664 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1666464484
transform 1 0 44620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1666464484
transform 1 0 48576 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1666464484
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1666464484
transform 1 0 56488 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1666464484
transform 1 0 3036 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1666464484
transform 1 0 6992 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1666464484
transform 1 0 10948 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1666464484
transform 1 0 14904 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1666464484
transform 1 0 18860 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1666464484
transform 1 0 22816 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1666464484
transform 1 0 26772 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1666464484
transform 1 0 30728 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1666464484
transform 1 0 34684 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1666464484
transform 1 0 38640 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1666464484
transform 1 0 42596 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1666464484
transform 1 0 46552 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1666464484
transform 1 0 50508 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1666464484
transform 1 0 54464 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1666464484
transform 1 0 58420 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1666464484
transform 1 0 5060 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1666464484
transform 1 0 9016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1666464484
transform 1 0 12972 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1666464484
transform 1 0 16928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1666464484
transform 1 0 20884 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1666464484
transform 1 0 24840 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1666464484
transform 1 0 28796 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1666464484
transform 1 0 32752 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1666464484
transform 1 0 36708 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1666464484
transform 1 0 40664 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1666464484
transform 1 0 44620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1666464484
transform 1 0 48576 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1666464484
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1666464484
transform 1 0 56488 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1666464484
transform 1 0 3036 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1666464484
transform 1 0 6992 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1666464484
transform 1 0 10948 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1666464484
transform 1 0 14904 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1666464484
transform 1 0 18860 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1666464484
transform 1 0 22816 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1666464484
transform 1 0 26772 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1666464484
transform 1 0 30728 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1666464484
transform 1 0 34684 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1666464484
transform 1 0 38640 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1666464484
transform 1 0 42596 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1666464484
transform 1 0 46552 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1666464484
transform 1 0 50508 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1666464484
transform 1 0 54464 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1666464484
transform 1 0 58420 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1666464484
transform 1 0 5060 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1666464484
transform 1 0 9016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1666464484
transform 1 0 12972 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1666464484
transform 1 0 16928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1666464484
transform 1 0 20884 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1666464484
transform 1 0 24840 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1666464484
transform 1 0 28796 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1666464484
transform 1 0 32752 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1666464484
transform 1 0 36708 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1666464484
transform 1 0 40664 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1666464484
transform 1 0 44620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1666464484
transform 1 0 48576 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1666464484
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1666464484
transform 1 0 56488 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1666464484
transform 1 0 3036 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1666464484
transform 1 0 6992 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1666464484
transform 1 0 10948 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1666464484
transform 1 0 14904 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1666464484
transform 1 0 18860 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1666464484
transform 1 0 22816 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1666464484
transform 1 0 26772 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1666464484
transform 1 0 30728 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1666464484
transform 1 0 34684 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1666464484
transform 1 0 38640 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1666464484
transform 1 0 42596 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1666464484
transform 1 0 46552 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1666464484
transform 1 0 50508 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1666464484
transform 1 0 54464 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1666464484
transform 1 0 58420 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1666464484
transform 1 0 5060 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1666464484
transform 1 0 9016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1666464484
transform 1 0 12972 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1666464484
transform 1 0 16928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1666464484
transform 1 0 20884 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1666464484
transform 1 0 24840 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1666464484
transform 1 0 28796 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1666464484
transform 1 0 32752 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1666464484
transform 1 0 36708 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1666464484
transform 1 0 40664 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1666464484
transform 1 0 44620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1666464484
transform 1 0 48576 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1666464484
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1666464484
transform 1 0 56488 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1666464484
transform 1 0 3036 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1666464484
transform 1 0 6992 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1666464484
transform 1 0 10948 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1666464484
transform 1 0 14904 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1666464484
transform 1 0 18860 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1666464484
transform 1 0 22816 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1666464484
transform 1 0 26772 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1666464484
transform 1 0 30728 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1666464484
transform 1 0 34684 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1666464484
transform 1 0 38640 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1666464484
transform 1 0 42596 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1666464484
transform 1 0 46552 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1666464484
transform 1 0 50508 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1666464484
transform 1 0 54464 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1666464484
transform 1 0 58420 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1666464484
transform 1 0 5060 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1666464484
transform 1 0 9016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1666464484
transform 1 0 12972 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1666464484
transform 1 0 16928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1666464484
transform 1 0 20884 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1666464484
transform 1 0 24840 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1666464484
transform 1 0 28796 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1666464484
transform 1 0 32752 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1666464484
transform 1 0 36708 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1666464484
transform 1 0 40664 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1666464484
transform 1 0 44620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1666464484
transform 1 0 48576 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1666464484
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1666464484
transform 1 0 56488 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1666464484
transform 1 0 3036 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1666464484
transform 1 0 6992 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1666464484
transform 1 0 10948 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1666464484
transform 1 0 14904 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1666464484
transform 1 0 18860 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1666464484
transform 1 0 22816 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1666464484
transform 1 0 26772 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1666464484
transform 1 0 30728 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1666464484
transform 1 0 34684 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1666464484
transform 1 0 38640 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1666464484
transform 1 0 42596 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1666464484
transform 1 0 46552 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1666464484
transform 1 0 50508 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1666464484
transform 1 0 54464 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1666464484
transform 1 0 58420 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1666464484
transform 1 0 5060 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1666464484
transform 1 0 9016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1666464484
transform 1 0 12972 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1666464484
transform 1 0 16928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1666464484
transform 1 0 20884 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1666464484
transform 1 0 24840 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1666464484
transform 1 0 28796 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1666464484
transform 1 0 32752 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1666464484
transform 1 0 36708 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1666464484
transform 1 0 40664 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1666464484
transform 1 0 44620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1666464484
transform 1 0 48576 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1666464484
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1666464484
transform 1 0 56488 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1666464484
transform 1 0 3036 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1666464484
transform 1 0 6992 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1666464484
transform 1 0 10948 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1666464484
transform 1 0 14904 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1666464484
transform 1 0 18860 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1666464484
transform 1 0 22816 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1666464484
transform 1 0 26772 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1666464484
transform 1 0 30728 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1666464484
transform 1 0 34684 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1666464484
transform 1 0 38640 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1666464484
transform 1 0 42596 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1666464484
transform 1 0 46552 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1666464484
transform 1 0 50508 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1666464484
transform 1 0 54464 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1666464484
transform 1 0 58420 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1666464484
transform 1 0 5060 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1666464484
transform 1 0 9016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1666464484
transform 1 0 12972 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1666464484
transform 1 0 16928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1666464484
transform 1 0 20884 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1666464484
transform 1 0 24840 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1666464484
transform 1 0 28796 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1666464484
transform 1 0 32752 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1666464484
transform 1 0 36708 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1666464484
transform 1 0 40664 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1666464484
transform 1 0 44620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1666464484
transform 1 0 48576 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1666464484
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1666464484
transform 1 0 56488 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1666464484
transform 1 0 3036 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1666464484
transform 1 0 6992 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1666464484
transform 1 0 10948 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1666464484
transform 1 0 14904 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1666464484
transform 1 0 18860 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1666464484
transform 1 0 22816 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1666464484
transform 1 0 26772 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1666464484
transform 1 0 30728 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1666464484
transform 1 0 34684 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1666464484
transform 1 0 38640 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1666464484
transform 1 0 42596 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1666464484
transform 1 0 46552 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1666464484
transform 1 0 50508 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1666464484
transform 1 0 54464 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1666464484
transform 1 0 58420 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1666464484
transform 1 0 5060 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1666464484
transform 1 0 9016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1666464484
transform 1 0 12972 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1666464484
transform 1 0 16928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1666464484
transform 1 0 20884 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1666464484
transform 1 0 24840 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1666464484
transform 1 0 28796 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1666464484
transform 1 0 32752 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1666464484
transform 1 0 36708 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1666464484
transform 1 0 40664 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1666464484
transform 1 0 44620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1666464484
transform 1 0 48576 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1666464484
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1666464484
transform 1 0 56488 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1666464484
transform 1 0 3036 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1666464484
transform 1 0 6992 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1666464484
transform 1 0 10948 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1666464484
transform 1 0 14904 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1666464484
transform 1 0 18860 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1666464484
transform 1 0 22816 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1666464484
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1666464484
transform 1 0 30728 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1666464484
transform 1 0 34684 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1666464484
transform 1 0 38640 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1666464484
transform 1 0 42596 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1666464484
transform 1 0 46552 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1666464484
transform 1 0 50508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1666464484
transform 1 0 54464 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1666464484
transform 1 0 58420 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1666464484
transform 1 0 5060 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1666464484
transform 1 0 9016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1666464484
transform 1 0 12972 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1666464484
transform 1 0 16928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1666464484
transform 1 0 20884 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1666464484
transform 1 0 24840 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1666464484
transform 1 0 28796 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1666464484
transform 1 0 32752 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1666464484
transform 1 0 36708 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1666464484
transform 1 0 40664 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1666464484
transform 1 0 44620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1666464484
transform 1 0 48576 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1666464484
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1666464484
transform 1 0 56488 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1666464484
transform 1 0 3036 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1666464484
transform 1 0 6992 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1666464484
transform 1 0 10948 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1666464484
transform 1 0 14904 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1666464484
transform 1 0 18860 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1666464484
transform 1 0 22816 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1666464484
transform 1 0 26772 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1666464484
transform 1 0 30728 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1666464484
transform 1 0 34684 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1666464484
transform 1 0 38640 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1666464484
transform 1 0 42596 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1666464484
transform 1 0 46552 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1666464484
transform 1 0 50508 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1666464484
transform 1 0 54464 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1666464484
transform 1 0 58420 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1666464484
transform 1 0 5060 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1666464484
transform 1 0 9016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1666464484
transform 1 0 12972 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1666464484
transform 1 0 16928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1666464484
transform 1 0 20884 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1666464484
transform 1 0 24840 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1666464484
transform 1 0 28796 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1666464484
transform 1 0 32752 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1666464484
transform 1 0 36708 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1666464484
transform 1 0 40664 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1666464484
transform 1 0 44620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1666464484
transform 1 0 48576 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1666464484
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1666464484
transform 1 0 56488 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1666464484
transform 1 0 3036 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1666464484
transform 1 0 6992 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1666464484
transform 1 0 10948 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1666464484
transform 1 0 14904 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1666464484
transform 1 0 18860 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1666464484
transform 1 0 22816 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1666464484
transform 1 0 26772 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1666464484
transform 1 0 30728 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1666464484
transform 1 0 34684 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1666464484
transform 1 0 38640 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1666464484
transform 1 0 42596 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1666464484
transform 1 0 46552 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1666464484
transform 1 0 50508 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1666464484
transform 1 0 54464 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1666464484
transform 1 0 58420 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1666464484
transform 1 0 5060 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1666464484
transform 1 0 9016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1666464484
transform 1 0 12972 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1666464484
transform 1 0 16928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1666464484
transform 1 0 20884 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1666464484
transform 1 0 24840 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1666464484
transform 1 0 28796 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1666464484
transform 1 0 32752 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1666464484
transform 1 0 36708 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1666464484
transform 1 0 40664 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1666464484
transform 1 0 44620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1666464484
transform 1 0 48576 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1666464484
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1666464484
transform 1 0 56488 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1666464484
transform 1 0 3036 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1666464484
transform 1 0 6992 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1666464484
transform 1 0 10948 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1666464484
transform 1 0 14904 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1666464484
transform 1 0 18860 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1666464484
transform 1 0 22816 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1666464484
transform 1 0 26772 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1666464484
transform 1 0 30728 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1666464484
transform 1 0 34684 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1666464484
transform 1 0 38640 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1666464484
transform 1 0 42596 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1666464484
transform 1 0 46552 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1666464484
transform 1 0 50508 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1666464484
transform 1 0 54464 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1666464484
transform 1 0 58420 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1666464484
transform 1 0 5060 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1666464484
transform 1 0 9016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1666464484
transform 1 0 12972 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1666464484
transform 1 0 16928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1666464484
transform 1 0 20884 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1666464484
transform 1 0 24840 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1666464484
transform 1 0 28796 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1666464484
transform 1 0 32752 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1666464484
transform 1 0 36708 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1666464484
transform 1 0 40664 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1666464484
transform 1 0 44620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1666464484
transform 1 0 48576 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1666464484
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1666464484
transform 1 0 56488 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1666464484
transform 1 0 3036 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1666464484
transform 1 0 6992 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1666464484
transform 1 0 10948 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1666464484
transform 1 0 14904 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1666464484
transform 1 0 18860 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1666464484
transform 1 0 22816 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1666464484
transform 1 0 26772 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1666464484
transform 1 0 30728 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1666464484
transform 1 0 34684 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1666464484
transform 1 0 38640 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1666464484
transform 1 0 42596 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1666464484
transform 1 0 46552 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1666464484
transform 1 0 50508 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1666464484
transform 1 0 54464 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1666464484
transform 1 0 58420 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1666464484
transform 1 0 5060 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1666464484
transform 1 0 9016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1666464484
transform 1 0 12972 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1666464484
transform 1 0 16928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1666464484
transform 1 0 20884 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1666464484
transform 1 0 24840 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1666464484
transform 1 0 28796 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1666464484
transform 1 0 32752 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1666464484
transform 1 0 36708 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1666464484
transform 1 0 40664 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1666464484
transform 1 0 44620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1666464484
transform 1 0 48576 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1666464484
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1666464484
transform 1 0 56488 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1666464484
transform 1 0 3036 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1666464484
transform 1 0 6992 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1666464484
transform 1 0 10948 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1666464484
transform 1 0 14904 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1666464484
transform 1 0 18860 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1666464484
transform 1 0 22816 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1666464484
transform 1 0 26772 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1666464484
transform 1 0 30728 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1666464484
transform 1 0 34684 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1666464484
transform 1 0 38640 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1666464484
transform 1 0 42596 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1666464484
transform 1 0 46552 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1666464484
transform 1 0 50508 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1666464484
transform 1 0 54464 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1666464484
transform 1 0 58420 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1666464484
transform 1 0 5060 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1666464484
transform 1 0 9016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1666464484
transform 1 0 12972 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1666464484
transform 1 0 16928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1666464484
transform 1 0 20884 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1666464484
transform 1 0 24840 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1666464484
transform 1 0 28796 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1666464484
transform 1 0 32752 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1666464484
transform 1 0 36708 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1666464484
transform 1 0 40664 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1666464484
transform 1 0 44620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1666464484
transform 1 0 48576 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1666464484
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1666464484
transform 1 0 56488 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1666464484
transform 1 0 3036 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1666464484
transform 1 0 6992 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1666464484
transform 1 0 10948 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1666464484
transform 1 0 14904 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1666464484
transform 1 0 18860 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1666464484
transform 1 0 22816 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1666464484
transform 1 0 26772 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1666464484
transform 1 0 30728 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1666464484
transform 1 0 34684 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1666464484
transform 1 0 38640 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1666464484
transform 1 0 42596 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1666464484
transform 1 0 46552 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1666464484
transform 1 0 50508 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1666464484
transform 1 0 54464 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1666464484
transform 1 0 58420 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1666464484
transform 1 0 5060 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1666464484
transform 1 0 9016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1666464484
transform 1 0 12972 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1666464484
transform 1 0 16928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1666464484
transform 1 0 20884 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1666464484
transform 1 0 24840 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1666464484
transform 1 0 28796 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1666464484
transform 1 0 32752 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1666464484
transform 1 0 36708 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1666464484
transform 1 0 40664 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1666464484
transform 1 0 44620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1666464484
transform 1 0 48576 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1666464484
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1666464484
transform 1 0 56488 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1666464484
transform 1 0 3036 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1666464484
transform 1 0 6992 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1666464484
transform 1 0 10948 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1666464484
transform 1 0 14904 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1666464484
transform 1 0 18860 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1666464484
transform 1 0 22816 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1666464484
transform 1 0 26772 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1666464484
transform 1 0 30728 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1666464484
transform 1 0 34684 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1666464484
transform 1 0 38640 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1666464484
transform 1 0 42596 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1666464484
transform 1 0 46552 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1666464484
transform 1 0 50508 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1666464484
transform 1 0 54464 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1666464484
transform 1 0 58420 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1666464484
transform 1 0 5060 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1666464484
transform 1 0 9016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1666464484
transform 1 0 12972 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1666464484
transform 1 0 16928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1666464484
transform 1 0 20884 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1666464484
transform 1 0 24840 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1666464484
transform 1 0 28796 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1666464484
transform 1 0 32752 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1666464484
transform 1 0 36708 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1666464484
transform 1 0 40664 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1666464484
transform 1 0 44620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1666464484
transform 1 0 48576 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1666464484
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1666464484
transform 1 0 56488 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1666464484
transform 1 0 3036 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1666464484
transform 1 0 6992 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1666464484
transform 1 0 10948 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1666464484
transform 1 0 14904 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1666464484
transform 1 0 18860 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1666464484
transform 1 0 22816 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1666464484
transform 1 0 26772 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1666464484
transform 1 0 30728 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1666464484
transform 1 0 34684 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1666464484
transform 1 0 38640 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1666464484
transform 1 0 42596 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1666464484
transform 1 0 46552 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1666464484
transform 1 0 50508 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1666464484
transform 1 0 54464 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1666464484
transform 1 0 58420 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1666464484
transform 1 0 5060 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1666464484
transform 1 0 9016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1666464484
transform 1 0 12972 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1666464484
transform 1 0 16928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1666464484
transform 1 0 20884 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1666464484
transform 1 0 24840 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1666464484
transform 1 0 28796 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1666464484
transform 1 0 32752 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1666464484
transform 1 0 36708 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1666464484
transform 1 0 40664 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1666464484
transform 1 0 44620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1666464484
transform 1 0 48576 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1666464484
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1666464484
transform 1 0 56488 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1666464484
transform 1 0 3036 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1666464484
transform 1 0 6992 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1666464484
transform 1 0 10948 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1666464484
transform 1 0 14904 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1666464484
transform 1 0 18860 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1666464484
transform 1 0 22816 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1666464484
transform 1 0 26772 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1666464484
transform 1 0 30728 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1666464484
transform 1 0 34684 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1666464484
transform 1 0 38640 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1666464484
transform 1 0 42596 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1666464484
transform 1 0 46552 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1666464484
transform 1 0 50508 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1666464484
transform 1 0 54464 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1666464484
transform 1 0 58420 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1666464484
transform 1 0 5060 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1666464484
transform 1 0 9016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1666464484
transform 1 0 12972 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1666464484
transform 1 0 16928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1666464484
transform 1 0 20884 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1666464484
transform 1 0 24840 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1666464484
transform 1 0 28796 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1666464484
transform 1 0 32752 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1666464484
transform 1 0 36708 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1666464484
transform 1 0 40664 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1666464484
transform 1 0 44620 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1666464484
transform 1 0 48576 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1666464484
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1666464484
transform 1 0 56488 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1666464484
transform 1 0 3036 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1666464484
transform 1 0 6992 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1666464484
transform 1 0 10948 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1666464484
transform 1 0 14904 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1666464484
transform 1 0 18860 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1666464484
transform 1 0 22816 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1666464484
transform 1 0 26772 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1666464484
transform 1 0 30728 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1666464484
transform 1 0 34684 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1666464484
transform 1 0 38640 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1666464484
transform 1 0 42596 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1666464484
transform 1 0 46552 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1666464484
transform 1 0 50508 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1666464484
transform 1 0 54464 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1666464484
transform 1 0 58420 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1666464484
transform 1 0 5060 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1666464484
transform 1 0 9016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1666464484
transform 1 0 12972 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1666464484
transform 1 0 16928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1666464484
transform 1 0 20884 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1666464484
transform 1 0 24840 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1666464484
transform 1 0 28796 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1666464484
transform 1 0 32752 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1666464484
transform 1 0 36708 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1666464484
transform 1 0 40664 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1666464484
transform 1 0 44620 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1666464484
transform 1 0 48576 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1666464484
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1666464484
transform 1 0 56488 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1666464484
transform 1 0 3036 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1666464484
transform 1 0 6992 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1666464484
transform 1 0 10948 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1666464484
transform 1 0 14904 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1666464484
transform 1 0 18860 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1666464484
transform 1 0 22816 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1666464484
transform 1 0 26772 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1666464484
transform 1 0 30728 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1666464484
transform 1 0 34684 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1666464484
transform 1 0 38640 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1666464484
transform 1 0 42596 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1666464484
transform 1 0 46552 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1666464484
transform 1 0 50508 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1666464484
transform 1 0 54464 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1666464484
transform 1 0 58420 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1666464484
transform 1 0 5060 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1666464484
transform 1 0 9016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1666464484
transform 1 0 12972 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1666464484
transform 1 0 16928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1666464484
transform 1 0 20884 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1666464484
transform 1 0 24840 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1666464484
transform 1 0 28796 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1666464484
transform 1 0 32752 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1666464484
transform 1 0 36708 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1666464484
transform 1 0 40664 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1666464484
transform 1 0 44620 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1666464484
transform 1 0 48576 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1666464484
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1666464484
transform 1 0 56488 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1666464484
transform 1 0 3036 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1666464484
transform 1 0 6992 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1666464484
transform 1 0 10948 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1666464484
transform 1 0 14904 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1666464484
transform 1 0 18860 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1666464484
transform 1 0 22816 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1666464484
transform 1 0 26772 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1666464484
transform 1 0 30728 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1666464484
transform 1 0 34684 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1666464484
transform 1 0 38640 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1666464484
transform 1 0 42596 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1666464484
transform 1 0 46552 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1666464484
transform 1 0 50508 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1666464484
transform 1 0 54464 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1666464484
transform 1 0 58420 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1666464484
transform 1 0 5060 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1666464484
transform 1 0 9016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1666464484
transform 1 0 12972 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1666464484
transform 1 0 16928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1666464484
transform 1 0 20884 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1666464484
transform 1 0 24840 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1666464484
transform 1 0 28796 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1666464484
transform 1 0 32752 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1666464484
transform 1 0 36708 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1666464484
transform 1 0 40664 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1666464484
transform 1 0 44620 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1666464484
transform 1 0 48576 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1666464484
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1666464484
transform 1 0 56488 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1666464484
transform 1 0 3036 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1666464484
transform 1 0 6992 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1666464484
transform 1 0 10948 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1666464484
transform 1 0 14904 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1666464484
transform 1 0 18860 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1666464484
transform 1 0 22816 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1666464484
transform 1 0 26772 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1666464484
transform 1 0 30728 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1666464484
transform 1 0 34684 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1666464484
transform 1 0 38640 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1666464484
transform 1 0 42596 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1666464484
transform 1 0 46552 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1666464484
transform 1 0 50508 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1666464484
transform 1 0 54464 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1666464484
transform 1 0 58420 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1666464484
transform 1 0 5060 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1666464484
transform 1 0 9016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1666464484
transform 1 0 12972 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1666464484
transform 1 0 16928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1666464484
transform 1 0 20884 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1666464484
transform 1 0 24840 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1666464484
transform 1 0 28796 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1666464484
transform 1 0 32752 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1666464484
transform 1 0 36708 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1666464484
transform 1 0 40664 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1666464484
transform 1 0 44620 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1666464484
transform 1 0 48576 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1666464484
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1666464484
transform 1 0 56488 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1666464484
transform 1 0 3036 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1666464484
transform 1 0 6992 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1666464484
transform 1 0 10948 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1666464484
transform 1 0 14904 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1666464484
transform 1 0 18860 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1666464484
transform 1 0 22816 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1666464484
transform 1 0 26772 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1666464484
transform 1 0 30728 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1666464484
transform 1 0 34684 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1666464484
transform 1 0 38640 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1666464484
transform 1 0 42596 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1666464484
transform 1 0 46552 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1666464484
transform 1 0 50508 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1666464484
transform 1 0 54464 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1666464484
transform 1 0 58420 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1666464484
transform 1 0 5060 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1666464484
transform 1 0 9016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1666464484
transform 1 0 12972 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1666464484
transform 1 0 16928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1666464484
transform 1 0 20884 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1666464484
transform 1 0 24840 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1666464484
transform 1 0 28796 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1666464484
transform 1 0 32752 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1666464484
transform 1 0 36708 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1666464484
transform 1 0 40664 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1666464484
transform 1 0 44620 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1666464484
transform 1 0 48576 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1666464484
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1666464484
transform 1 0 56488 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1666464484
transform 1 0 3036 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1666464484
transform 1 0 6992 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1666464484
transform 1 0 10948 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1666464484
transform 1 0 14904 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1666464484
transform 1 0 18860 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1666464484
transform 1 0 22816 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1666464484
transform 1 0 26772 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1666464484
transform 1 0 30728 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1666464484
transform 1 0 34684 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1666464484
transform 1 0 38640 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1666464484
transform 1 0 42596 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1666464484
transform 1 0 46552 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1666464484
transform 1 0 50508 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1666464484
transform 1 0 54464 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1666464484
transform 1 0 58420 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1666464484
transform 1 0 5060 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1666464484
transform 1 0 9016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1666464484
transform 1 0 12972 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1666464484
transform 1 0 16928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1666464484
transform 1 0 20884 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1666464484
transform 1 0 24840 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1666464484
transform 1 0 28796 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1666464484
transform 1 0 32752 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1666464484
transform 1 0 36708 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1666464484
transform 1 0 40664 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1666464484
transform 1 0 44620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1666464484
transform 1 0 48576 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1666464484
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1666464484
transform 1 0 56488 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1666464484
transform 1 0 3036 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1666464484
transform 1 0 6992 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1666464484
transform 1 0 10948 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1666464484
transform 1 0 14904 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1666464484
transform 1 0 18860 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1666464484
transform 1 0 22816 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1666464484
transform 1 0 26772 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1666464484
transform 1 0 30728 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1666464484
transform 1 0 34684 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1666464484
transform 1 0 38640 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1666464484
transform 1 0 42596 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1666464484
transform 1 0 46552 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1666464484
transform 1 0 50508 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1666464484
transform 1 0 54464 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1666464484
transform 1 0 58420 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1666464484
transform 1 0 5060 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1666464484
transform 1 0 9016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1666464484
transform 1 0 12972 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1666464484
transform 1 0 16928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1666464484
transform 1 0 20884 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1666464484
transform 1 0 24840 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1666464484
transform 1 0 28796 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1666464484
transform 1 0 32752 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1666464484
transform 1 0 36708 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1666464484
transform 1 0 40664 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1666464484
transform 1 0 44620 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1666464484
transform 1 0 48576 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1637
timestamp 1666464484
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1638
timestamp 1666464484
transform 1 0 56488 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1639
timestamp 1666464484
transform 1 0 3036 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1640
timestamp 1666464484
transform 1 0 6992 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1641
timestamp 1666464484
transform 1 0 10948 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1642
timestamp 1666464484
transform 1 0 14904 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1643
timestamp 1666464484
transform 1 0 18860 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1644
timestamp 1666464484
transform 1 0 22816 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1645
timestamp 1666464484
transform 1 0 26772 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1646
timestamp 1666464484
transform 1 0 30728 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1647
timestamp 1666464484
transform 1 0 34684 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1648
timestamp 1666464484
transform 1 0 38640 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1649
timestamp 1666464484
transform 1 0 42596 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1650
timestamp 1666464484
transform 1 0 46552 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1651
timestamp 1666464484
transform 1 0 50508 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1652
timestamp 1666464484
transform 1 0 54464 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1653
timestamp 1666464484
transform 1 0 58420 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1654
timestamp 1666464484
transform 1 0 5060 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1655
timestamp 1666464484
transform 1 0 9016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1656
timestamp 1666464484
transform 1 0 12972 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1657
timestamp 1666464484
transform 1 0 16928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1658
timestamp 1666464484
transform 1 0 20884 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1659
timestamp 1666464484
transform 1 0 24840 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1660
timestamp 1666464484
transform 1 0 28796 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1661
timestamp 1666464484
transform 1 0 32752 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1662
timestamp 1666464484
transform 1 0 36708 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1663
timestamp 1666464484
transform 1 0 40664 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1664
timestamp 1666464484
transform 1 0 44620 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1665
timestamp 1666464484
transform 1 0 48576 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1666
timestamp 1666464484
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1667
timestamp 1666464484
transform 1 0 56488 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1668
timestamp 1666464484
transform 1 0 3036 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1669
timestamp 1666464484
transform 1 0 6992 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1670
timestamp 1666464484
transform 1 0 10948 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1671
timestamp 1666464484
transform 1 0 14904 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1672
timestamp 1666464484
transform 1 0 18860 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1673
timestamp 1666464484
transform 1 0 22816 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1674
timestamp 1666464484
transform 1 0 26772 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1675
timestamp 1666464484
transform 1 0 30728 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1676
timestamp 1666464484
transform 1 0 34684 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1677
timestamp 1666464484
transform 1 0 38640 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1678
timestamp 1666464484
transform 1 0 42596 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1679
timestamp 1666464484
transform 1 0 46552 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1680
timestamp 1666464484
transform 1 0 50508 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1681
timestamp 1666464484
transform 1 0 54464 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1682
timestamp 1666464484
transform 1 0 58420 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1683
timestamp 1666464484
transform 1 0 3036 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1684
timestamp 1666464484
transform 1 0 4968 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1685
timestamp 1666464484
transform 1 0 6900 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1686
timestamp 1666464484
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1687
timestamp 1666464484
transform 1 0 10764 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1688
timestamp 1666464484
transform 1 0 12696 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1689
timestamp 1666464484
transform 1 0 14628 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1690
timestamp 1666464484
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1691
timestamp 1666464484
transform 1 0 18492 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1692
timestamp 1666464484
transform 1 0 20424 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1693
timestamp 1666464484
transform 1 0 22356 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1694
timestamp 1666464484
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1695
timestamp 1666464484
transform 1 0 26220 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1696
timestamp 1666464484
transform 1 0 28152 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1697
timestamp 1666464484
transform 1 0 30084 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1698
timestamp 1666464484
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1699
timestamp 1666464484
transform 1 0 33948 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1700
timestamp 1666464484
transform 1 0 35880 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1701
timestamp 1666464484
transform 1 0 37812 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1702
timestamp 1666464484
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1703
timestamp 1666464484
transform 1 0 41676 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1704
timestamp 1666464484
transform 1 0 43608 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1705
timestamp 1666464484
transform 1 0 45540 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1706
timestamp 1666464484
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1707
timestamp 1666464484
transform 1 0 49404 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1708
timestamp 1666464484
transform 1 0 51336 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1709
timestamp 1666464484
transform 1 0 53268 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1710
timestamp 1666464484
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1711
timestamp 1666464484
transform 1 0 57132 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _157_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26864 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _158_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26036 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _159_
timestamp 1666464484
transform 1 0 31004 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _160_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 38088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1666464484
transform 1 0 36800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1666464484
transform -1 0 37536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1666464484
transform 1 0 35328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1666464484
transform -1 0 35236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1666464484
transform -1 0 34224 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1666464484
transform 1 0 32108 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1666464484
transform -1 0 34408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1666464484
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1666464484
transform -1 0 34500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _170_
timestamp 1666464484
transform 1 0 29992 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1666464484
transform 1 0 31832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1666464484
transform 1 0 29348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1666464484
transform -1 0 29256 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1666464484
transform -1 0 31280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1666464484
transform 1 0 29992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1666464484
transform 1 0 29624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1666464484
transform -1 0 29624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1666464484
transform -1 0 27600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1666464484
transform -1 0 27968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1666464484
transform -1 0 27324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _181_
timestamp 1666464484
transform 1 0 25760 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1666464484
transform -1 0 25392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1666464484
transform 1 0 25760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1666464484
transform 1 0 27324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1666464484
transform 1 0 26036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1666464484
transform 1 0 23368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1666464484
transform -1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1666464484
transform -1 0 24104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1666464484
transform -1 0 21712 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1666464484
transform -1 0 24288 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1666464484
transform -1 0 26036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _193_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34500 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _194_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 35052 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _195_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 35604 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _196_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 28244 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _197_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34500 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _198_
timestamp 1666464484
transform -1 0 34132 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _199_
timestamp 1666464484
transform -1 0 30544 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _200_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 35512 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _201_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34408 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _202_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32660 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _203_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31924 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _204_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34040 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _205_
timestamp 1666464484
transform 1 0 32016 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _206_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29900 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _207_
timestamp 1666464484
transform -1 0 30544 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _208_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29256 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _209_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35420 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _210_
timestamp 1666464484
transform -1 0 27416 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _211_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28612 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _212_
timestamp 1666464484
transform 1 0 28060 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _213_
timestamp 1666464484
transform -1 0 45356 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _214_
timestamp 1666464484
transform 1 0 43240 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _215_
timestamp 1666464484
transform -1 0 43516 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _216_
timestamp 1666464484
transform -1 0 38640 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _217_
timestamp 1666464484
transform 1 0 43884 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _218_
timestamp 1666464484
transform -1 0 43516 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _219_
timestamp 1666464484
transform -1 0 39376 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _220_
timestamp 1666464484
transform -1 0 42320 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _221_
timestamp 1666464484
transform -1 0 42504 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _222_
timestamp 1666464484
transform -1 0 42320 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _223_
timestamp 1666464484
transform -1 0 40480 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _224_
timestamp 1666464484
transform -1 0 41400 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _225_
timestamp 1666464484
transform 1 0 40388 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _226_
timestamp 1666464484
transform -1 0 38456 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _227_
timestamp 1666464484
transform -1 0 39376 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _228_
timestamp 1666464484
transform 1 0 37812 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _229_
timestamp 1666464484
transform 1 0 44252 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _230_
timestamp 1666464484
transform 1 0 37168 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _231_
timestamp 1666464484
transform 1 0 37812 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _232_
timestamp 1666464484
transform -1 0 35604 0 1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _233_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 36156 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _234_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27968 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _235_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28152 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1666464484
transform -1 0 35696 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _237_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31648 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _238_
timestamp 1666464484
transform 1 0 31188 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _239_
timestamp 1666464484
transform 1 0 30728 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1666464484
transform -1 0 39836 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _241_
timestamp 1666464484
transform -1 0 41216 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _242_
timestamp 1666464484
transform 1 0 40940 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _243_
timestamp 1666464484
transform 1 0 40020 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _244_
timestamp 1666464484
transform -1 0 25024 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _245_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22356 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _246_
timestamp 1666464484
transform -1 0 24472 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1666464484
transform -1 0 23644 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _248_
timestamp 1666464484
transform -1 0 24380 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _249_
timestamp 1666464484
transform -1 0 33580 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _250_
timestamp 1666464484
transform 1 0 32108 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _251_
timestamp 1666464484
transform 1 0 33948 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _252_
timestamp 1666464484
transform 1 0 33212 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _253_
timestamp 1666464484
transform 1 0 33028 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _254_
timestamp 1666464484
transform -1 0 41860 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _255_
timestamp 1666464484
transform 1 0 40756 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _256_
timestamp 1666464484
transform 1 0 42872 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _257_
timestamp 1666464484
transform 1 0 41584 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _258_
timestamp 1666464484
transform 1 0 41860 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _259_
timestamp 1666464484
transform -1 0 25852 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1666464484
transform 1 0 25300 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _261_
timestamp 1666464484
transform -1 0 25668 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1666464484
transform -1 0 24840 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _263_
timestamp 1666464484
transform -1 0 25760 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _264_
timestamp 1666464484
transform 1 0 32108 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _265_
timestamp 1666464484
transform 1 0 30084 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _266_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31648 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _267_
timestamp 1666464484
transform 1 0 30912 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _268_
timestamp 1666464484
transform -1 0 31280 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _269_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31004 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _270_
timestamp 1666464484
transform 1 0 43884 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _271_
timestamp 1666464484
transform -1 0 41492 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _272_
timestamp 1666464484
transform 1 0 38824 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _273_
timestamp 1666464484
transform 1 0 39744 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _274_
timestamp 1666464484
transform -1 0 39836 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _275_
timestamp 1666464484
transform 1 0 39560 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _276_
timestamp 1666464484
transform -1 0 26588 0 1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1666464484
transform 1 0 25944 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _278_
timestamp 1666464484
transform -1 0 27416 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _279_
timestamp 1666464484
transform -1 0 26864 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _280_
timestamp 1666464484
transform -1 0 27784 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _281_
timestamp 1666464484
transform 1 0 29348 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _282_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28060 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _283_
timestamp 1666464484
transform 1 0 28796 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _284_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29256 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _285_
timestamp 1666464484
transform 1 0 32016 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _286_
timestamp 1666464484
transform 1 0 33028 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _287_
timestamp 1666464484
transform -1 0 28428 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _288_
timestamp 1666464484
transform 1 0 37904 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _289_
timestamp 1666464484
transform -1 0 38548 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _290_
timestamp 1666464484
transform -1 0 37628 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _291_
timestamp 1666464484
transform 1 0 43884 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _292_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 43884 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _293_
timestamp 1666464484
transform 1 0 36340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _294_
timestamp 1666464484
transform 1 0 35972 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _295_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29164 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _296_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28888 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _519__194 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 25668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24656 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _520_
timestamp 1666464484
transform 1 0 22724 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _520__195
timestamp 1666464484
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _521_
timestamp 1666464484
transform 1 0 25760 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _521__196
timestamp 1666464484
transform 1 0 22356 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _522_
timestamp 1666464484
transform -1 0 22632 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _522__197
timestamp 1666464484
transform 1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _523_
timestamp 1666464484
transform 1 0 22724 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _523__198
timestamp 1666464484
transform -1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _524__199
timestamp 1666464484
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _524_
timestamp 1666464484
transform 1 0 24656 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _525_
timestamp 1666464484
transform 1 0 26680 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _525__200
timestamp 1666464484
transform 1 0 26036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _526_
timestamp 1666464484
transform 1 0 27508 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _526__201
timestamp 1666464484
transform 1 0 27324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _527__202
timestamp 1666464484
transform -1 0 28336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _527_
timestamp 1666464484
transform 1 0 26680 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _528_
timestamp 1666464484
transform 1 0 27968 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _528__203
timestamp 1666464484
transform 1 0 25392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _529__204
timestamp 1666464484
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _529_
timestamp 1666464484
transform -1 0 24656 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _530_
timestamp 1666464484
transform -1 0 26588 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _530__205
timestamp 1666464484
transform 1 0 25392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _531_
timestamp 1666464484
transform 1 0 26680 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _531__206
timestamp 1666464484
transform 1 0 26036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _532_
timestamp 1666464484
transform 1 0 26680 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _532__207
timestamp 1666464484
transform -1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _533__208
timestamp 1666464484
transform 1 0 27968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _533_
timestamp 1666464484
transform 1 0 28612 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _534__209
timestamp 1666464484
transform -1 0 30544 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _534_
timestamp 1666464484
transform 1 0 29532 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _535__210
timestamp 1666464484
transform 1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _535_
timestamp 1666464484
transform 1 0 30084 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _536_
timestamp 1666464484
transform 1 0 30084 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _536__211
timestamp 1666464484
transform -1 0 30636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _537_
timestamp 1666464484
transform 1 0 28612 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _537__212
timestamp 1666464484
transform -1 0 29900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _538_
timestamp 1666464484
transform 1 0 30636 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _538__213
timestamp 1666464484
transform -1 0 31280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _539__214
timestamp 1666464484
transform -1 0 31280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _539_
timestamp 1666464484
transform 1 0 31004 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _540_
timestamp 1666464484
transform -1 0 34960 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _540__215
timestamp 1666464484
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _541_
timestamp 1666464484
transform 1 0 34960 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _541__216
timestamp 1666464484
transform -1 0 35604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _542_
timestamp 1666464484
transform -1 0 33764 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _542__217
timestamp 1666464484
transform 1 0 32292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _543__218
timestamp 1666464484
transform -1 0 33580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _543_
timestamp 1666464484
transform 1 0 32016 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _544__219
timestamp 1666464484
transform -1 0 33304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _544_
timestamp 1666464484
transform 1 0 33028 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _545__220
timestamp 1666464484
transform -1 0 35696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _545_
timestamp 1666464484
transform -1 0 35052 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _546_
timestamp 1666464484
transform 1 0 36984 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _546__221
timestamp 1666464484
transform 1 0 35972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _547_
timestamp 1666464484
transform -1 0 36892 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _547__222
timestamp 1666464484
transform 1 0 35972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _548_
timestamp 1666464484
transform 1 0 36984 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _548__223
timestamp 1666464484
transform 1 0 36156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _549_
timestamp 1666464484
transform -1 0 35880 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _549__224
timestamp 1666464484
transform -1 0 38180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _550__225
timestamp 1666464484
transform 1 0 34960 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _550_
timestamp 1666464484
transform -1 0 36156 0 -1 53312
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3772 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform -1 0 28612 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform -1 0 30544 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1666464484
transform 1 0 35880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1666464484
transform 1 0 34592 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1666464484
transform 1 0 36156 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1666464484
transform 1 0 38088 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1666464484
transform 1 0 38916 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1666464484
transform -1 0 41216 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1666464484
transform 1 0 46552 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1666464484
transform -1 0 43424 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1666464484
transform 1 0 44896 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1666464484
transform -1 0 46184 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1666464484
transform 1 0 47748 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1666464484
transform 1 0 48392 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1666464484
transform 1 0 49772 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 51612 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 53084 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1666464484
transform 1 0 53912 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1666464484
transform 1 0 55476 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  macro_10_37
timestamp 1666464484
transform -1 0 51060 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_38
timestamp 1666464484
transform -1 0 52348 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_39
timestamp 1666464484
transform -1 0 53636 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_40
timestamp 1666464484
transform -1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_41
timestamp 1666464484
transform -1 0 56488 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_42
timestamp 1666464484
transform -1 0 6716 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_43
timestamp 1666464484
transform -1 0 8004 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_44
timestamp 1666464484
transform -1 0 9568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_45
timestamp 1666464484
transform -1 0 30268 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_46
timestamp 1666464484
transform -1 0 34500 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_47
timestamp 1666464484
transform -1 0 36432 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_48
timestamp 1666464484
transform -1 0 36800 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_49
timestamp 1666464484
transform -1 0 37444 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_50
timestamp 1666464484
transform -1 0 40020 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_51
timestamp 1666464484
transform -1 0 39192 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_52
timestamp 1666464484
transform -1 0 40480 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_53
timestamp 1666464484
transform -1 0 46092 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_54
timestamp 1666464484
transform -1 0 45264 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_55
timestamp 1666464484
transform -1 0 47104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_56
timestamp 1666464484
transform -1 0 45908 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_57
timestamp 1666464484
transform -1 0 47288 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_58
timestamp 1666464484
transform -1 0 49956 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_59
timestamp 1666464484
transform -1 0 49772 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_60
timestamp 1666464484
transform -1 0 51704 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_61
timestamp 1666464484
transform -1 0 52992 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_62
timestamp 1666464484
transform -1 0 54280 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_63
timestamp 1666464484
transform -1 0 55108 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_64
timestamp 1666464484
transform -1 0 56488 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_65
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_66
timestamp 1666464484
transform -1 0 17940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_67
timestamp 1666464484
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_68
timestamp 1666464484
transform 1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_69
timestamp 1666464484
transform -1 0 18768 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_70
timestamp 1666464484
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_71
timestamp 1666464484
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_72
timestamp 1666464484
transform -1 0 19596 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_73
timestamp 1666464484
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_74
timestamp 1666464484
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_75
timestamp 1666464484
transform 1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_76
timestamp 1666464484
transform -1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_77
timestamp 1666464484
transform 1 0 19780 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_78
timestamp 1666464484
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_79
timestamp 1666464484
transform 1 0 18492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_80
timestamp 1666464484
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_81
timestamp 1666464484
transform 1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_82
timestamp 1666464484
transform 1 0 20424 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_83
timestamp 1666464484
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_84
timestamp 1666464484
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_85
timestamp 1666464484
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_86
timestamp 1666464484
transform -1 0 23460 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_87
timestamp 1666464484
transform 1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_88
timestamp 1666464484
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_89
timestamp 1666464484
transform -1 0 24288 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_90
timestamp 1666464484
transform 1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_91
timestamp 1666464484
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_92
timestamp 1666464484
transform 1 0 19320 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_93
timestamp 1666464484
transform 1 0 20424 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_94
timestamp 1666464484
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_95
timestamp 1666464484
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_96
timestamp 1666464484
transform 1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_97
timestamp 1666464484
transform -1 0 39008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_98
timestamp 1666464484
transform -1 0 36340 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_99
timestamp 1666464484
transform -1 0 40296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_100
timestamp 1666464484
transform -1 0 39560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_101
timestamp 1666464484
transform -1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_102
timestamp 1666464484
transform -1 0 37536 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_103
timestamp 1666464484
transform -1 0 39192 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_104
timestamp 1666464484
transform -1 0 40204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_105
timestamp 1666464484
transform -1 0 38180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_106
timestamp 1666464484
transform -1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_107
timestamp 1666464484
transform -1 0 39560 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_108
timestamp 1666464484
transform -1 0 39192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_109
timestamp 1666464484
transform -1 0 41216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_110
timestamp 1666464484
transform -1 0 40480 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_111
timestamp 1666464484
transform -1 0 42228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_112
timestamp 1666464484
transform -1 0 40204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_113
timestamp 1666464484
transform -1 0 41124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_114
timestamp 1666464484
transform -1 0 41860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_115
timestamp 1666464484
transform -1 0 42872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_116
timestamp 1666464484
transform -1 0 41216 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_117
timestamp 1666464484
transform -1 0 42504 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_118
timestamp 1666464484
transform -1 0 41768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_119
timestamp 1666464484
transform -1 0 43148 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_120
timestamp 1666464484
transform -1 0 42412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_121
timestamp 1666464484
transform -1 0 44160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_122
timestamp 1666464484
transform -1 0 43792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_123
timestamp 1666464484
transform -1 0 43148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_124
timestamp 1666464484
transform -1 0 44804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_125
timestamp 1666464484
transform -1 0 43792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_126
timestamp 1666464484
transform -1 0 44436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_127
timestamp 1666464484
transform -1 0 44436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_128
timestamp 1666464484
transform -1 0 45172 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_129
timestamp 1666464484
transform -1 0 46092 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_130
timestamp 1666464484
transform -1 0 45080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_131
timestamp 1666464484
transform -1 0 45816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_132
timestamp 1666464484
transform -1 0 46736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_133
timestamp 1666464484
transform -1 0 45724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_134
timestamp 1666464484
transform -1 0 46460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_135
timestamp 1666464484
transform -1 0 46368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_136
timestamp 1666464484
transform -1 0 47104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_137
timestamp 1666464484
transform -1 0 48024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_138
timestamp 1666464484
transform -1 0 47104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_139
timestamp 1666464484
transform -1 0 47748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_140
timestamp 1666464484
transform -1 0 48668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_141
timestamp 1666464484
transform -1 0 47748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_142
timestamp 1666464484
transform -1 0 48392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_143
timestamp 1666464484
transform -1 0 48392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_144
timestamp 1666464484
transform -1 0 49128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_145
timestamp 1666464484
transform -1 0 49956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_146
timestamp 1666464484
transform -1 0 50600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_147
timestamp 1666464484
transform -1 0 49772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_148
timestamp 1666464484
transform -1 0 49404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_149
timestamp 1666464484
transform -1 0 50416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_150
timestamp 1666464484
transform -1 0 50048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_151
timestamp 1666464484
transform -1 0 51060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_152
timestamp 1666464484
transform -1 0 51888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_153
timestamp 1666464484
transform -1 0 52532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_154
timestamp 1666464484
transform -1 0 51704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_155
timestamp 1666464484
transform -1 0 51336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_156
timestamp 1666464484
transform -1 0 52348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_157
timestamp 1666464484
transform -1 0 51980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_158
timestamp 1666464484
transform -1 0 53820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_159
timestamp 1666464484
transform -1 0 53084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_160
timestamp 1666464484
transform -1 0 54464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_161
timestamp 1666464484
transform 1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_162
timestamp 1666464484
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_163
timestamp 1666464484
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_164
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_165
timestamp 1666464484
transform -1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_166
timestamp 1666464484
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_167
timestamp 1666464484
transform 1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_168
timestamp 1666464484
transform -1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_169
timestamp 1666464484
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_170
timestamp 1666464484
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_171
timestamp 1666464484
transform 1 0 10580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_172
timestamp 1666464484
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_173
timestamp 1666464484
transform 1 0 11224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_174
timestamp 1666464484
transform -1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_175
timestamp 1666464484
transform 1 0 11868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_176
timestamp 1666464484
transform 1 0 11592 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_177
timestamp 1666464484
transform -1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_178
timestamp 1666464484
transform 1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_179
timestamp 1666464484
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_180
timestamp 1666464484
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_181
timestamp 1666464484
transform 1 0 13248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_182
timestamp 1666464484
transform 1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_183
timestamp 1666464484
transform -1 0 14720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_184
timestamp 1666464484
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_185
timestamp 1666464484
transform -1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_186
timestamp 1666464484
transform 1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_187
timestamp 1666464484
transform 1 0 14168 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_188
timestamp 1666464484
transform -1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_189
timestamp 1666464484
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_190
timestamp 1666464484
transform -1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_191
timestamp 1666464484
transform 1 0 15824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_192
timestamp 1666464484
transform 1 0 16468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_193
timestamp 1666464484
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_226
timestamp 1666464484
transform -1 0 4784 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_227
timestamp 1666464484
transform -1 0 6348 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_228
timestamp 1666464484
transform -1 0 7728 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_229
timestamp 1666464484
transform 1 0 8372 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_230
timestamp 1666464484
transform -1 0 10488 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_231
timestamp 1666464484
transform -1 0 11868 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_232
timestamp 1666464484
transform -1 0 13248 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_233
timestamp 1666464484
transform -1 0 14444 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_234
timestamp 1666464484
transform -1 0 16008 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_235
timestamp 1666464484
transform -1 0 17388 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_236
timestamp 1666464484
transform -1 0 19412 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_237
timestamp 1666464484
transform -1 0 20148 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_238
timestamp 1666464484
transform -1 0 21528 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_239
timestamp 1666464484
transform -1 0 22908 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_240
timestamp 1666464484
transform -1 0 24196 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_241
timestamp 1666464484
transform -1 0 25668 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_242
timestamp 1666464484
transform 1 0 25208 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_243
timestamp 1666464484
transform 1 0 27508 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_244
timestamp 1666464484
transform -1 0 29808 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_245
timestamp 1666464484
transform -1 0 31280 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_246
timestamp 1666464484
transform -1 0 35604 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_247
timestamp 1666464484
transform -1 0 39192 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_248
timestamp 1666464484
transform -1 0 36340 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_249
timestamp 1666464484
transform -1 0 37260 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_250
timestamp 1666464484
transform -1 0 38088 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_251
timestamp 1666464484
transform -1 0 45080 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_252
timestamp 1666464484
transform -1 0 45448 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_253
timestamp 1666464484
transform -1 0 43148 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_254
timestamp 1666464484
transform -1 0 46000 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_255
timestamp 1666464484
transform -1 0 46644 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_256
timestamp 1666464484
transform -1 0 47748 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_257
timestamp 1666464484
transform -1 0 47932 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_10_258
timestamp 1666464484
transform -1 0 49128 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1666464484
transform -1 0 5612 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1666464484
transform -1 0 19320 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1666464484
transform -1 0 21068 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1666464484
transform -1 0 22080 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1666464484
transform -1 0 23368 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1666464484
transform 1 0 23736 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1666464484
transform 1 0 25852 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1666464484
transform 1 0 27232 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1666464484
transform 1 0 30360 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1666464484
transform -1 0 11408 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1666464484
transform -1 0 12420 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1666464484
transform -1 0 13800 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1666464484
transform -1 0 15272 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1666464484
transform -1 0 17204 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1666464484
transform -1 0 17940 0 -1 57664
box -38 -48 406 592
<< labels >>
flabel metal2 s 3698 59200 3754 60000 0 FreeSans 224 90 0 0 io_active
port 0 nsew signal input
flabel metal2 s 4158 59200 4214 60000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 17958 59200 18014 60000 0 FreeSans 224 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s 19338 59200 19394 60000 0 FreeSans 224 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal2 s 20718 59200 20774 60000 0 FreeSans 224 90 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 22098 59200 22154 60000 0 FreeSans 224 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 23478 59200 23534 60000 0 FreeSans 224 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal2 s 24858 59200 24914 60000 0 FreeSans 224 90 0 0 io_in[15]
port 7 nsew signal input
flabel metal2 s 26238 59200 26294 60000 0 FreeSans 224 90 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 27618 59200 27674 60000 0 FreeSans 224 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 28998 59200 29054 60000 0 FreeSans 224 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 30378 59200 30434 60000 0 FreeSans 224 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal2 s 5538 59200 5594 60000 0 FreeSans 224 90 0 0 io_in[1]
port 12 nsew signal input
flabel metal2 s 31758 59200 31814 60000 0 FreeSans 224 90 0 0 io_in[20]
port 13 nsew signal input
flabel metal2 s 33138 59200 33194 60000 0 FreeSans 224 90 0 0 io_in[21]
port 14 nsew signal input
flabel metal2 s 34518 59200 34574 60000 0 FreeSans 224 90 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 35898 59200 35954 60000 0 FreeSans 224 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 37278 59200 37334 60000 0 FreeSans 224 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 38658 59200 38714 60000 0 FreeSans 224 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 40038 59200 40094 60000 0 FreeSans 224 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal2 s 41418 59200 41474 60000 0 FreeSans 224 90 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 42798 59200 42854 60000 0 FreeSans 224 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 44178 59200 44234 60000 0 FreeSans 224 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 6918 59200 6974 60000 0 FreeSans 224 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal2 s 45558 59200 45614 60000 0 FreeSans 224 90 0 0 io_in[30]
port 24 nsew signal input
flabel metal2 s 46938 59200 46994 60000 0 FreeSans 224 90 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 48318 59200 48374 60000 0 FreeSans 224 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal2 s 49698 59200 49754 60000 0 FreeSans 224 90 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 51078 59200 51134 60000 0 FreeSans 224 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 52458 59200 52514 60000 0 FreeSans 224 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal2 s 53838 59200 53894 60000 0 FreeSans 224 90 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 55218 59200 55274 60000 0 FreeSans 224 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 8298 59200 8354 60000 0 FreeSans 224 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal2 s 9678 59200 9734 60000 0 FreeSans 224 90 0 0 io_in[4]
port 33 nsew signal input
flabel metal2 s 11058 59200 11114 60000 0 FreeSans 224 90 0 0 io_in[5]
port 34 nsew signal input
flabel metal2 s 12438 59200 12494 60000 0 FreeSans 224 90 0 0 io_in[6]
port 35 nsew signal input
flabel metal2 s 13818 59200 13874 60000 0 FreeSans 224 90 0 0 io_in[7]
port 36 nsew signal input
flabel metal2 s 15198 59200 15254 60000 0 FreeSans 224 90 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 16578 59200 16634 60000 0 FreeSans 224 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 4618 59200 4674 60000 0 FreeSans 224 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal2 s 18418 59200 18474 60000 0 FreeSans 224 90 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal2 s 19798 59200 19854 60000 0 FreeSans 224 90 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal2 s 21178 59200 21234 60000 0 FreeSans 224 90 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal2 s 22558 59200 22614 60000 0 FreeSans 224 90 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal2 s 23938 59200 23994 60000 0 FreeSans 224 90 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 25318 59200 25374 60000 0 FreeSans 224 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal2 s 26698 59200 26754 60000 0 FreeSans 224 90 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 28078 59200 28134 60000 0 FreeSans 224 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 29458 59200 29514 60000 0 FreeSans 224 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 30838 59200 30894 60000 0 FreeSans 224 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal2 s 5998 59200 6054 60000 0 FreeSans 224 90 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal2 s 32218 59200 32274 60000 0 FreeSans 224 90 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal2 s 33598 59200 33654 60000 0 FreeSans 224 90 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 34978 59200 35034 60000 0 FreeSans 224 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 36358 59200 36414 60000 0 FreeSans 224 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 37738 59200 37794 60000 0 FreeSans 224 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal2 s 39118 59200 39174 60000 0 FreeSans 224 90 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal2 s 40498 59200 40554 60000 0 FreeSans 224 90 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 41878 59200 41934 60000 0 FreeSans 224 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal2 s 43258 59200 43314 60000 0 FreeSans 224 90 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal2 s 44638 59200 44694 60000 0 FreeSans 224 90 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 7378 59200 7434 60000 0 FreeSans 224 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal2 s 46018 59200 46074 60000 0 FreeSans 224 90 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal2 s 47398 59200 47454 60000 0 FreeSans 224 90 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal2 s 48778 59200 48834 60000 0 FreeSans 224 90 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal2 s 50158 59200 50214 60000 0 FreeSans 224 90 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal2 s 51538 59200 51594 60000 0 FreeSans 224 90 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal2 s 52918 59200 52974 60000 0 FreeSans 224 90 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal2 s 54298 59200 54354 60000 0 FreeSans 224 90 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal2 s 55678 59200 55734 60000 0 FreeSans 224 90 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 8758 59200 8814 60000 0 FreeSans 224 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal2 s 10138 59200 10194 60000 0 FreeSans 224 90 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal2 s 11518 59200 11574 60000 0 FreeSans 224 90 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal2 s 12898 59200 12954 60000 0 FreeSans 224 90 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 14278 59200 14334 60000 0 FreeSans 224 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 15658 59200 15714 60000 0 FreeSans 224 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 17038 59200 17094 60000 0 FreeSans 224 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal2 s 5078 59200 5134 60000 0 FreeSans 224 90 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal2 s 18878 59200 18934 60000 0 FreeSans 224 90 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal2 s 20258 59200 20314 60000 0 FreeSans 224 90 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal2 s 21638 59200 21694 60000 0 FreeSans 224 90 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal2 s 23018 59200 23074 60000 0 FreeSans 224 90 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal2 s 24398 59200 24454 60000 0 FreeSans 224 90 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal2 s 25778 59200 25834 60000 0 FreeSans 224 90 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal2 s 27158 59200 27214 60000 0 FreeSans 224 90 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 28538 59200 28594 60000 0 FreeSans 224 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal2 s 29918 59200 29974 60000 0 FreeSans 224 90 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal2 s 31298 59200 31354 60000 0 FreeSans 224 90 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 6458 59200 6514 60000 0 FreeSans 224 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 32678 59200 32734 60000 0 FreeSans 224 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal2 s 34058 59200 34114 60000 0 FreeSans 224 90 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 35438 59200 35494 60000 0 FreeSans 224 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal2 s 36818 59200 36874 60000 0 FreeSans 224 90 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 38198 59200 38254 60000 0 FreeSans 224 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 39578 59200 39634 60000 0 FreeSans 224 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal2 s 40958 59200 41014 60000 0 FreeSans 224 90 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 42338 59200 42394 60000 0 FreeSans 224 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 43718 59200 43774 60000 0 FreeSans 224 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal2 s 45098 59200 45154 60000 0 FreeSans 224 90 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 7838 59200 7894 60000 0 FreeSans 224 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal2 s 46478 59200 46534 60000 0 FreeSans 224 90 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal2 s 47858 59200 47914 60000 0 FreeSans 224 90 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal2 s 49238 59200 49294 60000 0 FreeSans 224 90 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal2 s 50618 59200 50674 60000 0 FreeSans 224 90 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal2 s 51998 59200 52054 60000 0 FreeSans 224 90 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal2 s 53378 59200 53434 60000 0 FreeSans 224 90 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 54758 59200 54814 60000 0 FreeSans 224 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal2 s 56138 59200 56194 60000 0 FreeSans 224 90 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal2 s 9218 59200 9274 60000 0 FreeSans 224 90 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal2 s 10598 59200 10654 60000 0 FreeSans 224 90 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 11978 59200 12034 60000 0 FreeSans 224 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 13358 59200 13414 60000 0 FreeSans 224 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal2 s 14738 59200 14794 60000 0 FreeSans 224 90 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 16118 59200 16174 60000 0 FreeSans 224 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal2 s 17498 59200 17554 60000 0 FreeSans 224 90 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 115 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 116 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 117 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 118 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 119 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 120 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 121 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 122 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 123 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 124 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 125 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 126 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 127 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 128 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 129 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 130 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 131 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 132 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 133 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 134 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 135 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 136 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 137 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 138 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 139 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 140 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 141 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 142 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 143 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 144 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 145 nsew signal input
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 146 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 147 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 148 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 149 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 150 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 151 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 152 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 153 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 154 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 155 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 156 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 157 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 158 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 159 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 160 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 161 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 162 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 163 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 164 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 165 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 166 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 167 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 168 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 169 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 170 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 171 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 172 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 173 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 174 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 175 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 176 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 177 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 178 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 179 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 180 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 181 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 182 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 183 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 184 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 185 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 186 nsew signal input
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 187 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 188 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 189 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 190 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 191 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 192 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 193 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 194 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 195 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 196 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 197 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 198 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 199 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 200 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 201 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 202 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 203 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 204 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 205 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 206 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 207 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 208 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 209 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 210 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 211 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 212 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 213 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 214 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 215 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 216 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 217 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 218 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 219 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 220 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 221 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 222 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 223 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 224 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 225 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 226 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 227 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 228 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 229 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 230 nsew signal input
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 231 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 232 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 233 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 234 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 235 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 236 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 237 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 238 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 239 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 240 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 241 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 242 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 243 nsew signal tristate
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 244 nsew signal tristate
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 245 nsew signal tristate
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 246 nsew signal tristate
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 247 nsew signal tristate
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 248 nsew signal tristate
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 249 nsew signal tristate
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 250 nsew signal tristate
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 251 nsew signal tristate
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 252 nsew signal tristate
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 253 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 254 nsew signal tristate
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 255 nsew signal tristate
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 256 nsew signal tristate
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 257 nsew signal tristate
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 258 nsew signal tristate
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 259 nsew signal tristate
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 260 nsew signal tristate
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 261 nsew signal tristate
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 262 nsew signal tristate
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 263 nsew signal tristate
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 264 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 265 nsew signal tristate
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 266 nsew signal tristate
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 267 nsew signal tristate
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 268 nsew signal tristate
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 269 nsew signal tristate
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 270 nsew signal tristate
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 271 nsew signal tristate
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 272 nsew signal tristate
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 273 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 274 nsew signal tristate
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 275 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 276 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 277 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 278 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 279 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 280 nsew signal tristate
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 281 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 282 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 283 nsew signal tristate
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 284 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 285 nsew signal tristate
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 286 nsew signal tristate
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 287 nsew signal tristate
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 288 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 289 nsew signal tristate
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 290 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 291 nsew signal tristate
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 292 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 293 nsew signal tristate
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 294 nsew signal tristate
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 295 nsew signal tristate
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 296 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 297 nsew signal tristate
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 298 nsew signal tristate
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 299 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 300 nsew signal tristate
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 301 nsew signal tristate
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 302 nsew signal tristate
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 303 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 304 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 305 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 306 nsew signal tristate
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 307 nsew signal tristate
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 308 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 309 nsew signal tristate
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 310 nsew signal tristate
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 311 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 312 nsew signal tristate
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 313 nsew signal tristate
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 314 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 315 nsew signal tristate
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 316 nsew signal tristate
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 317 nsew signal tristate
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 318 nsew signal tristate
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 319 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 320 nsew signal tristate
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 321 nsew signal tristate
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 322 nsew signal tristate
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 323 nsew signal tristate
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 324 nsew signal tristate
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 325 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 326 nsew signal tristate
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 327 nsew signal tristate
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 328 nsew signal tristate
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 329 nsew signal tristate
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 330 nsew signal tristate
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 331 nsew signal tristate
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 332 nsew signal tristate
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 333 nsew signal tristate
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 334 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 335 nsew signal tristate
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 336 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 337 nsew signal tristate
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 338 nsew signal tristate
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 339 nsew signal tristate
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 340 nsew signal tristate
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 341 nsew signal tristate
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 342 nsew signal tristate
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 343 nsew signal tristate
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 344 nsew signal tristate
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 345 nsew signal tristate
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 346 nsew signal tristate
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 347 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 348 nsew signal tristate
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 349 nsew signal tristate
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 350 nsew signal tristate
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 351 nsew signal tristate
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 352 nsew signal tristate
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 353 nsew signal tristate
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 354 nsew signal tristate
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 355 nsew signal tristate
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 356 nsew signal tristate
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 357 nsew signal tristate
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 358 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 359 nsew signal tristate
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 360 nsew signal tristate
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 361 nsew signal tristate
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 362 nsew signal tristate
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 363 nsew signal tristate
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 364 nsew signal tristate
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 365 nsew signal tristate
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 366 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 367 nsew signal tristate
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 368 nsew signal tristate
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 369 nsew signal tristate
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 370 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 371 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 372 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 373 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 374 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 375 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 376 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 377 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 378 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 379 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 380 nsew signal input
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 381 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 382 nsew signal input
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 383 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 384 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 385 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 386 nsew signal input
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 387 nsew signal input
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 388 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 389 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 390 nsew signal input
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 391 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 392 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 393 nsew signal input
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 394 nsew signal input
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 395 nsew signal input
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 396 nsew signal input
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 397 nsew signal input
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 398 nsew signal input
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 399 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 400 nsew signal input
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 401 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 402 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 403 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 404 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 405 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 406 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 407 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 408 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 409 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 410 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 411 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 412 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 413 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 414 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 415 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 416 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 417 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 418 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 419 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 420 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 421 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 422 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 423 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 424 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 425 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 426 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 427 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 428 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 429 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 430 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 431 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 432 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 433 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 434 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 435 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 436 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 437 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 438 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 439 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 440 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 441 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 442 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 443 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 444 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 445 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 446 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 447 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 448 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 449 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 450 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 451 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 452 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 453 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 454 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 455 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 456 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 457 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 458 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 459 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 460 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 461 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 462 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 463 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 464 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 465 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 466 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 467 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 468 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 469 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 470 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 471 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 472 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 473 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 474 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 475 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 476 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 477 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 478 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 479 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 480 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 481 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 482 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 483 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 484 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 485 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 486 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 487 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 488 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 489 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 490 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 491 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 492 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 493 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 494 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 495 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 496 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 497 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 498 nsew signal input
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 500 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 500 nsew ground bidirectional
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wb_clk_i
port 501 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wb_rst_i
port 502 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 503 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 504 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 505 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 506 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 507 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 508 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 509 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 510 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 511 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 512 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 513 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 514 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 515 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 516 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 517 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 518 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 519 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 520 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 521 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 522 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 523 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 524 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 525 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 526 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 527 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 528 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 529 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 530 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 531 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 532 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 533 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 534 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 535 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 536 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 537 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 538 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 539 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 540 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 541 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 542 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 543 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 544 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 545 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 546 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 547 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 548 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 549 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 550 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 551 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 552 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 553 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 554 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 555 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 556 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 557 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 558 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 559 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 560 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 561 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 562 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 563 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 564 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 565 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 566 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 567 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 568 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 569 nsew signal tristate
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 570 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 571 nsew signal tristate
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 572 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 573 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 574 nsew signal tristate
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 575 nsew signal tristate
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 576 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 577 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 578 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 579 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 580 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 581 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 582 nsew signal tristate
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 583 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 584 nsew signal tristate
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 585 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 586 nsew signal tristate
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 587 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 588 nsew signal tristate
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 589 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 590 nsew signal tristate
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 591 nsew signal tristate
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 592 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 593 nsew signal tristate
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 594 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 595 nsew signal tristate
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 596 nsew signal tristate
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 597 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 598 nsew signal tristate
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 599 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 600 nsew signal tristate
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 601 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 602 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 603 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 604 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 605 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_we_i
port 606 nsew signal input
rlabel metal1 29992 57120 29992 57120 0 vccd1
rlabel metal1 29992 57664 29992 57664 0 vssd1
rlabel metal2 34546 55420 34546 55420 0 _000_
rlabel metal2 35512 55318 35512 55318 0 _001_
rlabel metal1 29348 56338 29348 56338 0 _002_
rlabel metal1 28704 55114 28704 55114 0 _003_
rlabel metal1 34270 54094 34270 54094 0 _004_
rlabel metal2 33534 54434 33534 54434 0 _005_
rlabel metal2 29578 54774 29578 54774 0 _006_
rlabel metal1 34132 53754 34132 53754 0 _007_
rlabel metal2 33166 54026 33166 54026 0 _008_
rlabel metal1 32614 54298 32614 54298 0 _009_
rlabel metal2 32430 54876 32430 54876 0 _010_
rlabel metal1 33534 55046 33534 55046 0 _011_
rlabel metal1 30958 54128 30958 54128 0 _012_
rlabel metal1 29762 55284 29762 55284 0 _013_
rlabel metal1 30084 54502 30084 54502 0 _014_
rlabel metal1 28060 55726 28060 55726 0 _015_
rlabel metal1 27370 55624 27370 55624 0 _016_
rlabel metal2 28290 56168 28290 56168 0 _017_
rlabel metal1 28014 56406 28014 56406 0 _018_
rlabel metal1 28612 56474 28612 56474 0 _019_
rlabel metal1 41860 55182 41860 55182 0 _020_
rlabel metal1 43792 55658 43792 55658 0 _021_
rlabel metal1 38226 54706 38226 54706 0 _022_
rlabel metal2 37398 54774 37398 54774 0 _023_
rlabel metal1 43654 55182 43654 55182 0 _024_
rlabel metal1 38962 55148 38962 55148 0 _025_
rlabel metal1 38134 55692 38134 55692 0 _026_
rlabel metal2 41906 54842 41906 54842 0 _027_
rlabel metal2 41814 55012 41814 55012 0 _028_
rlabel metal1 41906 55726 41906 55726 0 _029_
rlabel metal2 40894 55216 40894 55216 0 _030_
rlabel metal1 40618 55760 40618 55760 0 _031_
rlabel metal2 39790 55080 39790 55080 0 _032_
rlabel metal1 38272 55726 38272 55726 0 _033_
rlabel metal1 38134 55284 38134 55284 0 _034_
rlabel metal1 37950 55930 37950 55930 0 _035_
rlabel metal1 38318 56882 38318 56882 0 _036_
rlabel metal2 35834 55862 35834 55862 0 _037_
rlabel metal1 35558 56848 35558 56848 0 _038_
rlabel metal1 34960 57018 34960 57018 0 _039_
rlabel metal2 33718 55556 33718 55556 0 _040_
rlabel metal1 31556 57018 31556 57018 0 _041_
rlabel metal1 31234 56202 31234 56202 0 _042_
rlabel metal1 24242 56270 24242 56270 0 _043_
rlabel metal2 36754 56304 36754 56304 0 _044_
rlabel metal2 41170 56508 41170 56508 0 _045_
rlabel metal1 40756 56474 40756 56474 0 _046_
rlabel metal2 40066 57698 40066 57698 0 _047_
rlabel metal1 22632 56814 22632 56814 0 _048_
rlabel metal1 23736 56338 23736 56338 0 _049_
rlabel metal1 32706 54638 32706 54638 0 _050_
rlabel metal1 33074 54774 33074 54774 0 _051_
rlabel metal1 33902 56474 33902 56474 0 _052_
rlabel metal2 33258 56508 33258 56508 0 _053_
rlabel metal1 25438 56406 25438 56406 0 _054_
rlabel metal2 40986 55114 40986 55114 0 _055_
rlabel metal2 42274 55318 42274 55318 0 _056_
rlabel metal1 42555 56814 42555 56814 0 _057_
rlabel metal1 42044 56338 42044 56338 0 _058_
rlabel metal1 25622 56678 25622 56678 0 _059_
rlabel metal2 25530 56236 25530 56236 0 _060_
rlabel metal2 24610 55930 24610 55930 0 _061_
rlabel metal1 31326 55624 31326 55624 0 _062_
rlabel metal1 31188 55736 31188 55736 0 _063_
rlabel metal1 31096 54842 31096 54842 0 _064_
rlabel metal1 31418 55386 31418 55386 0 _065_
rlabel metal1 31464 54026 31464 54026 0 _066_
rlabel metal1 27186 56270 27186 56270 0 _067_
rlabel metal1 41906 56406 41906 56406 0 _068_
rlabel metal1 39790 56406 39790 56406 0 _069_
rlabel metal2 39606 54672 39606 54672 0 _070_
rlabel metal2 40158 55590 40158 55590 0 _071_
rlabel metal1 39790 54060 39790 54060 0 _072_
rlabel metal1 39560 56474 39560 56474 0 _073_
rlabel metal2 26174 55964 26174 55964 0 _074_
rlabel metal2 26634 55692 26634 55692 0 _075_
rlabel metal2 29394 54332 29394 54332 0 _076_
rlabel metal2 29118 55046 29118 55046 0 _077_
rlabel metal1 29532 54774 29532 54774 0 _078_
rlabel metal1 29256 53754 29256 53754 0 _079_
rlabel metal1 29348 56814 29348 56814 0 _080_
rlabel metal2 28566 55760 28566 55760 0 _081_
rlabel metal2 28382 56032 28382 56032 0 _082_
rlabel metal2 37950 55862 37950 55862 0 _083_
rlabel metal1 37766 56270 37766 56270 0 _084_
rlabel metal1 36938 56474 36938 56474 0 _085_
rlabel metal2 43930 57052 43930 57052 0 _086_
rlabel metal2 36294 56882 36294 56882 0 _087_
rlabel metal1 36248 55794 36248 55794 0 _088_
rlabel metal2 26082 5440 26082 5440 0 _089_
rlabel metal1 37490 2414 37490 2414 0 _090_
rlabel metal2 30314 5984 30314 5984 0 _091_
rlabel metal1 23414 2380 23414 2380 0 _092_
rlabel metal2 24886 6188 24886 6188 0 _093_
rlabel metal1 23552 5270 23552 5270 0 _094_
rlabel metal1 23276 3162 23276 3162 0 _095_
rlabel metal1 23920 2618 23920 2618 0 _096_
rlabel metal1 23138 2618 23138 2618 0 _097_
rlabel metal1 24196 4522 24196 4522 0 _098_
rlabel metal1 26542 6358 26542 6358 0 _099_
rlabel metal2 27002 5474 27002 5474 0 _100_
rlabel metal2 26910 5950 26910 5950 0 _101_
rlabel metal2 28198 4522 28198 4522 0 _102_
rlabel metal2 25254 2788 25254 2788 0 _103_
rlabel metal1 26772 2618 26772 2618 0 _104_
rlabel metal2 27830 2788 27830 2788 0 _105_
rlabel metal2 27462 3876 27462 3876 0 _106_
rlabel metal2 29486 3842 29486 3842 0 _107_
rlabel metal2 29762 6766 29762 6766 0 _108_
rlabel metal1 30222 4250 30222 4250 0 _109_
rlabel metal2 31142 2788 31142 2788 0 _110_
rlabel metal2 29118 3026 29118 3026 0 _111_
rlabel metal1 30866 4012 30866 4012 0 _112_
rlabel metal2 31234 5916 31234 5916 0 _113_
rlabel metal1 34546 2618 34546 2618 0 _114_
rlabel metal1 35190 2618 35190 2618 0 _115_
rlabel metal1 33902 3434 33902 3434 0 _116_
rlabel metal2 32246 5644 32246 5644 0 _117_
rlabel metal2 33258 4794 33258 4794 0 _118_
rlabel metal2 34822 5406 34822 5406 0 _119_
rlabel metal2 35466 3502 35466 3502 0 _120_
rlabel metal2 37398 4114 37398 4114 0 _121_
rlabel metal1 37076 2550 37076 2550 0 _122_
rlabel metal2 38226 4488 38226 4488 0 _123_
rlabel metal2 36018 57358 36018 57358 0 _124_
rlabel metal1 3818 57494 3818 57494 0 io_active
rlabel metal1 28704 54162 28704 54162 0 io_in[18]
rlabel metal1 30406 55250 30406 55250 0 io_in[19]
rlabel metal1 34914 57426 34914 57426 0 io_in[20]
rlabel metal1 36018 54638 36018 54638 0 io_in[21]
rlabel metal1 37444 57494 37444 57494 0 io_in[22]
rlabel metal2 36202 55012 36202 55012 0 io_in[23]
rlabel metal1 37720 57358 37720 57358 0 io_in[24]
rlabel metal1 38824 56882 38824 56882 0 io_in[25]
rlabel metal1 40664 54162 40664 54162 0 io_in[26]
rlabel metal1 44252 55590 44252 55590 0 io_in[27]
rlabel metal1 43102 57426 43102 57426 0 io_in[28]
rlabel metal1 44666 55250 44666 55250 0 io_in[29]
rlabel metal1 45816 57426 45816 57426 0 io_in[30]
rlabel metal1 47380 57426 47380 57426 0 io_in[31]
rlabel metal1 48392 56882 48392 56882 0 io_in[32]
rlabel metal1 49772 57426 49772 57426 0 io_in[33]
rlabel metal1 51382 57426 51382 57426 0 io_in[34]
rlabel metal1 52716 57494 52716 57494 0 io_in[35]
rlabel metal1 53912 57426 53912 57426 0 io_in[36]
rlabel metal1 55384 57426 55384 57426 0 io_in[37]
rlabel metal1 5244 57562 5244 57562 0 io_out[0]
rlabel metal1 18998 57562 18998 57562 0 io_out[10]
rlabel metal1 20562 57562 20562 57562 0 io_out[11]
rlabel metal1 21758 57562 21758 57562 0 io_out[12]
rlabel metal1 23092 57562 23092 57562 0 io_out[13]
rlabel metal1 24196 57562 24196 57562 0 io_out[14]
rlabel metal1 25944 55930 25944 55930 0 io_out[15]
rlabel metal1 27370 55386 27370 55386 0 io_out[16]
rlabel metal1 29946 57290 29946 57290 0 io_out[17]
rlabel metal1 11132 57562 11132 57562 0 io_out[4]
rlabel metal1 12098 57562 12098 57562 0 io_out[5]
rlabel metal1 13478 57562 13478 57562 0 io_out[6]
rlabel metal1 14904 57562 14904 57562 0 io_out[7]
rlabel metal2 16146 58388 16146 58388 0 io_out[8]
rlabel metal1 17618 57562 17618 57562 0 io_out[9]
rlabel metal2 26174 3254 26174 3254 0 la_data_out[32]
rlabel metal2 25438 3978 25438 3978 0 la_data_out[33]
rlabel metal2 26726 2115 26726 2115 0 la_data_out[34]
rlabel metal1 22034 3604 22034 3604 0 la_data_out[35]
rlabel metal1 25415 4046 25415 4046 0 la_data_out[36]
rlabel metal2 27554 2642 27554 2642 0 la_data_out[37]
rlabel metal2 27830 1639 27830 1639 0 la_data_out[38]
rlabel metal2 28106 3254 28106 3254 0 la_data_out[39]
rlabel metal2 28382 2948 28382 2948 0 la_data_out[40]
rlabel metal2 28658 3798 28658 3798 0 la_data_out[41]
rlabel metal1 24150 2924 24150 2924 0 la_data_out[42]
rlabel metal2 29210 2200 29210 2200 0 la_data_out[43]
rlabel metal2 29486 1860 29486 1860 0 la_data_out[44]
rlabel metal2 29762 2404 29762 2404 0 la_data_out[45]
rlabel metal2 30038 2710 30038 2710 0 la_data_out[46]
rlabel metal2 30314 1979 30314 1979 0 la_data_out[47]
rlabel metal2 30590 2948 30590 2948 0 la_data_out[48]
rlabel metal2 30866 1826 30866 1826 0 la_data_out[49]
rlabel metal2 31142 1231 31142 1231 0 la_data_out[50]
rlabel metal2 31418 2404 31418 2404 0 la_data_out[51]
rlabel metal2 31694 3254 31694 3254 0 la_data_out[52]
rlabel metal2 31970 1860 31970 1860 0 la_data_out[53]
rlabel metal2 32246 2200 32246 2200 0 la_data_out[54]
rlabel metal2 32522 2166 32522 2166 0 la_data_out[55]
rlabel metal2 32798 2710 32798 2710 0 la_data_out[56]
rlabel metal2 33074 2370 33074 2370 0 la_data_out[57]
rlabel metal2 33350 2948 33350 2948 0 la_data_out[58]
rlabel metal1 36110 2958 36110 2958 0 la_data_out[59]
rlabel metal2 33902 2336 33902 2336 0 la_data_out[60]
rlabel metal1 37490 3978 37490 3978 0 la_data_out[61]
rlabel metal2 34454 3492 34454 3492 0 la_data_out[62]
rlabel metal2 34730 1639 34730 1639 0 la_data_out[63]
rlabel metal2 16974 56984 16974 56984 0 net1
rlabel metal1 40388 55046 40388 55046 0 net10
rlabel metal1 36018 2856 36018 2856 0 net100
rlabel metal2 36110 1554 36110 1554 0 net101
rlabel metal2 36386 1962 36386 1962 0 net102
rlabel metal2 36662 2200 36662 2200 0 net103
rlabel metal2 36938 2098 36938 2098 0 net104
rlabel metal2 37214 1571 37214 1571 0 net105
rlabel metal2 37490 1299 37490 1299 0 net106
rlabel metal2 37766 2336 37766 2336 0 net107
rlabel metal2 38042 1826 38042 1826 0 net108
rlabel metal2 38318 1095 38318 1095 0 net109
rlabel metal1 43148 56814 43148 56814 0 net11
rlabel metal2 38594 2166 38594 2166 0 net110
rlabel metal2 38870 1622 38870 1622 0 net111
rlabel metal2 39146 2370 39146 2370 0 net112
rlabel metal2 39422 2200 39422 2200 0 net113
rlabel metal2 39698 1860 39698 1860 0 net114
rlabel metal2 39974 1656 39974 1656 0 net115
rlabel metal2 40250 2336 40250 2336 0 net116
rlabel metal2 40526 1826 40526 1826 0 net117
rlabel metal2 40802 2166 40802 2166 0 net118
rlabel metal2 41078 1894 41078 1894 0 net119
rlabel metal1 39146 55692 39146 55692 0 net12
rlabel metal2 41354 2132 41354 2132 0 net120
rlabel metal2 41630 1554 41630 1554 0 net121
rlabel metal2 41906 1860 41906 1860 0 net122
rlabel metal2 42182 2200 42182 2200 0 net123
rlabel metal2 42458 1622 42458 1622 0 net124
rlabel metal2 42734 2132 42734 2132 0 net125
rlabel metal2 43010 1826 43010 1826 0 net126
rlabel metal2 43286 2200 43286 2200 0 net127
rlabel metal2 43562 1792 43562 1792 0 net128
rlabel metal2 43838 1656 43838 1656 0 net129
rlabel metal1 39238 54706 39238 54706 0 net13
rlabel metal2 44114 2166 44114 2166 0 net130
rlabel metal2 44390 1860 44390 1860 0 net131
rlabel metal2 44666 1622 44666 1622 0 net132
rlabel metal2 44942 2132 44942 2132 0 net133
rlabel metal2 45218 1826 45218 1826 0 net134
rlabel metal2 45494 2200 45494 2200 0 net135
rlabel metal2 45770 1792 45770 1792 0 net136
rlabel metal2 46046 1588 46046 1588 0 net137
rlabel metal2 46322 2132 46322 2132 0 net138
rlabel metal2 46598 1860 46598 1860 0 net139
rlabel metal1 45172 55182 45172 55182 0 net14
rlabel metal2 46874 1656 46874 1656 0 net140
rlabel metal2 47150 2132 47150 2132 0 net141
rlabel metal2 47426 1826 47426 1826 0 net142
rlabel metal2 47702 2132 47702 2132 0 net143
rlabel metal2 47978 1792 47978 1792 0 net144
rlabel metal2 48254 1622 48254 1622 0 net145
rlabel metal2 48530 1588 48530 1588 0 net146
rlabel metal2 48806 1826 48806 1826 0 net147
rlabel metal2 49082 2132 49082 2132 0 net148
rlabel metal2 49358 1792 49358 1792 0 net149
rlabel metal2 43378 57188 43378 57188 0 net15
rlabel metal2 49634 2132 49634 2132 0 net150
rlabel metal2 49910 1860 49910 1860 0 net151
rlabel metal2 50186 1622 50186 1622 0 net152
rlabel metal2 50462 1027 50462 1027 0 net153
rlabel metal2 50738 1826 50738 1826 0 net154
rlabel metal2 51014 2132 51014 2132 0 net155
rlabel metal2 51290 1792 51290 1792 0 net156
rlabel metal2 51566 2132 51566 2132 0 net157
rlabel metal2 51842 1656 51842 1656 0 net158
rlabel metal2 52118 1860 52118 1860 0 net159
rlabel metal2 44114 56287 44114 56287 0 net16
rlabel metal2 52394 1622 52394 1622 0 net160
rlabel metal2 7682 1792 7682 1792 0 net161
rlabel metal2 8234 1792 8234 1792 0 net162
rlabel metal2 8602 1656 8602 1656 0 net163
rlabel metal2 8970 1792 8970 1792 0 net164
rlabel metal2 9338 2132 9338 2132 0 net165
rlabel metal2 9706 1588 9706 1588 0 net166
rlabel metal2 9982 1792 9982 1792 0 net167
rlabel metal2 10258 2132 10258 2132 0 net168
rlabel metal2 10534 1792 10534 1792 0 net169
rlabel metal1 47242 57358 47242 57358 0 net17
rlabel metal2 10810 1622 10810 1622 0 net170
rlabel metal2 11086 1792 11086 1792 0 net171
rlabel metal2 11362 1588 11362 1588 0 net172
rlabel metal2 11638 1792 11638 1792 0 net173
rlabel metal2 11914 2132 11914 2132 0 net174
rlabel metal2 12190 1792 12190 1792 0 net175
rlabel metal2 12466 1656 12466 1656 0 net176
rlabel metal2 12742 2132 12742 2132 0 net177
rlabel metal2 13018 1792 13018 1792 0 net178
rlabel metal2 13294 1588 13294 1588 0 net179
rlabel metal1 39836 57426 39836 57426 0 net18
rlabel metal2 13570 2132 13570 2132 0 net180
rlabel metal2 13846 1792 13846 1792 0 net181
rlabel metal2 14122 1792 14122 1792 0 net182
rlabel metal2 14398 2132 14398 2132 0 net183
rlabel metal2 14674 1622 14674 1622 0 net184
rlabel metal2 14950 2132 14950 2132 0 net185
rlabel metal2 15226 1792 15226 1792 0 net186
rlabel metal2 15502 1588 15502 1588 0 net187
rlabel metal2 15778 2132 15778 2132 0 net188
rlabel metal2 16054 1860 16054 1860 0 net189
rlabel metal2 40434 57630 40434 57630 0 net19
rlabel metal2 16330 2336 16330 2336 0 net190
rlabel metal2 16606 1792 16606 1792 0 net191
rlabel metal2 16882 2132 16882 2132 0 net192
rlabel metal2 17158 1622 17158 1622 0 net193
rlabel metal2 24702 5916 24702 5916 0 net194
rlabel metal2 22310 4624 22310 4624 0 net195
rlabel metal1 24196 7310 24196 7310 0 net196
rlabel metal1 22448 3026 22448 3026 0 net197
rlabel metal1 23092 3706 23092 3706 0 net198
rlabel metal1 24472 4590 24472 4590 0 net199
rlabel metal2 32062 54502 32062 54502 0 net2
rlabel metal2 54142 56984 54142 56984 0 net20
rlabel metal2 26266 5168 26266 5168 0 net200
rlabel metal2 27554 5236 27554 5236 0 net201
rlabel metal1 27416 7174 27416 7174 0 net202
rlabel metal2 25622 5474 25622 5474 0 net203
rlabel metal2 24610 3264 24610 3264 0 net204
rlabel metal2 26542 3264 26542 3264 0 net205
rlabel metal1 26496 2958 26496 2958 0 net206
rlabel metal2 28014 3842 28014 3842 0 net207
rlabel metal1 28428 4590 28428 4590 0 net208
rlabel metal2 29578 6528 29578 6528 0 net209
rlabel metal2 54234 56304 54234 56304 0 net21
rlabel metal1 29900 5134 29900 5134 0 net210
rlabel metal2 30406 2754 30406 2754 0 net211
rlabel metal2 29670 3094 29670 3094 0 net212
rlabel metal1 30866 3706 30866 3706 0 net213
rlabel metal2 31050 6256 31050 6256 0 net214
rlabel metal1 33856 2550 33856 2550 0 net215
rlabel metal1 35190 3026 35190 3026 0 net216
rlabel metal1 33120 2618 33120 2618 0 net217
rlabel metal1 32062 4692 32062 4692 0 net218
rlabel metal2 33074 5100 33074 5100 0 net219
rlabel metal1 5566 57392 5566 57392 0 net22
rlabel metal1 35236 5134 35236 5134 0 net220
rlabel metal1 36202 2992 36202 2992 0 net221
rlabel metal1 36524 4114 36524 4114 0 net222
rlabel metal1 36708 2618 36708 2618 0 net223
rlabel metal2 37950 4964 37950 4964 0 net224
rlabel metal2 36110 53312 36110 53312 0 net225
rlabel metal1 4600 57426 4600 57426 0 net226
rlabel metal1 6072 57018 6072 57018 0 net227
rlabel metal1 7452 57018 7452 57018 0 net228
rlabel metal1 8694 57426 8694 57426 0 net229
rlabel metal2 19274 57188 19274 57188 0 net23
rlabel metal1 10212 57426 10212 57426 0 net230
rlabel metal1 11592 57018 11592 57018 0 net231
rlabel metal1 12972 57018 12972 57018 0 net232
rlabel metal1 14260 57426 14260 57426 0 net233
rlabel metal1 15732 57426 15732 57426 0 net234
rlabel metal1 17112 57018 17112 57018 0 net235
rlabel metal1 18814 57018 18814 57018 0 net236
rlabel metal1 19964 57426 19964 57426 0 net237
rlabel metal1 21252 57018 21252 57018 0 net238
rlabel metal1 22632 56338 22632 56338 0 net239
rlabel metal2 21022 57596 21022 57596 0 net24
rlabel metal2 23966 57572 23966 57572 0 net240
rlabel metal1 25392 54842 25392 54842 0 net241
rlabel metal1 26082 55862 26082 55862 0 net242
rlabel metal1 27922 54842 27922 54842 0 net243
rlabel metal1 29532 53074 29532 53074 0 net244
rlabel metal1 30958 57018 30958 57018 0 net245
rlabel metal2 35374 56814 35374 56814 0 net246
rlabel metal1 37628 56134 37628 56134 0 net247
rlabel metal2 36110 54876 36110 54876 0 net248
rlabel metal1 36708 54162 36708 54162 0 net249
rlabel metal2 22034 57630 22034 57630 0 net25
rlabel metal1 37812 53754 37812 53754 0 net250
rlabel metal2 39146 57861 39146 57861 0 net251
rlabel metal2 40618 56916 40618 56916 0 net252
rlabel metal2 42918 55658 42918 55658 0 net253
rlabel metal1 44528 56202 44528 56202 0 net254
rlabel metal1 45540 56270 45540 56270 0 net255
rlabel metal1 46782 57018 46782 57018 0 net256
rlabel metal1 47564 56338 47564 56338 0 net257
rlabel metal1 48852 56338 48852 56338 0 net258
rlabel metal1 23322 57460 23322 57460 0 net26
rlabel metal2 23782 56644 23782 56644 0 net27
rlabel metal1 24978 55930 24978 55930 0 net28
rlabel metal1 27140 55250 27140 55250 0 net29
rlabel metal1 32154 53550 32154 53550 0 net3
rlabel metal1 30406 57392 30406 57392 0 net30
rlabel metal2 21390 57086 21390 57086 0 net31
rlabel via2 12374 57443 12374 57443 0 net32
rlabel metal1 13754 57460 13754 57460 0 net33
rlabel metal2 15226 57664 15226 57664 0 net34
rlabel metal1 17158 57324 17158 57324 0 net35
rlabel metal1 17894 57392 17894 57392 0 net36
rlabel metal1 50508 57018 50508 57018 0 net37
rlabel metal1 51842 57018 51842 57018 0 net38
rlabel metal1 53176 57018 53176 57018 0 net39
rlabel metal2 32614 56542 32614 56542 0 net4
rlabel metal1 54510 57426 54510 57426 0 net40
rlabel metal1 55982 57426 55982 57426 0 net41
rlabel metal2 6486 58320 6486 58320 0 net42
rlabel metal1 7820 57426 7820 57426 0 net43
rlabel metal1 9292 57426 9292 57426 0 net44
rlabel metal1 29992 53754 29992 53754 0 net45
rlabel metal2 34270 57290 34270 57290 0 net46
rlabel metal1 36110 55182 36110 55182 0 net47
rlabel metal2 36570 55352 36570 55352 0 net48
rlabel metal2 37214 55386 37214 55386 0 net49
rlabel metal2 28014 55964 28014 55964 0 net5
rlabel metal1 38364 55862 38364 55862 0 net50
rlabel metal1 38916 53754 38916 53754 0 net51
rlabel metal1 40158 53958 40158 53958 0 net52
rlabel metal2 41078 56763 41078 56763 0 net53
rlabel metal1 44896 55930 44896 55930 0 net54
rlabel metal1 45310 56950 45310 56950 0 net55
rlabel metal1 45402 55930 45402 55930 0 net56
rlabel metal1 46782 56338 46782 56338 0 net57
rlabel metal1 48806 57018 48806 57018 0 net58
rlabel metal1 49404 56338 49404 56338 0 net59
rlabel metal1 31756 56814 31756 56814 0 net6
rlabel metal2 50646 58082 50646 58082 0 net60
rlabel metal1 52624 57018 52624 57018 0 net61
rlabel metal1 53774 57018 53774 57018 0 net62
rlabel metal1 54832 57018 54832 57018 0 net63
rlabel metal1 56212 57018 56212 57018 0 net64
rlabel metal2 17342 1792 17342 1792 0 net65
rlabel metal2 17618 2336 17618 2336 0 net66
rlabel metal2 17894 2132 17894 2132 0 net67
rlabel metal2 18170 2132 18170 2132 0 net68
rlabel metal2 18446 2336 18446 2336 0 net69
rlabel metal2 34454 56814 34454 56814 0 net7
rlabel metal2 18722 1656 18722 1656 0 net70
rlabel metal2 18998 1860 18998 1860 0 net71
rlabel metal2 19274 1775 19274 1775 0 net72
rlabel metal2 19550 1095 19550 1095 0 net73
rlabel metal2 19826 1367 19826 1367 0 net74
rlabel metal2 20102 2166 20102 2166 0 net75
rlabel metal2 20378 2676 20378 2676 0 net76
rlabel metal2 20654 2404 20654 2404 0 net77
rlabel metal2 20930 1622 20930 1622 0 net78
rlabel metal2 21206 1894 21206 1894 0 net79
rlabel metal1 35190 55250 35190 55250 0 net8
rlabel metal2 21482 2200 21482 2200 0 net80
rlabel metal2 21758 2676 21758 2676 0 net81
rlabel metal2 22034 2370 22034 2370 0 net82
rlabel metal2 22310 1554 22310 1554 0 net83
rlabel metal2 22586 1826 22586 1826 0 net84
rlabel metal2 22862 2880 22862 2880 0 net85
rlabel metal2 23138 3220 23138 3220 0 net86
rlabel metal2 23414 2744 23414 2744 0 net87
rlabel metal2 23690 2064 23690 2064 0 net88
rlabel metal2 23966 3424 23966 3424 0 net89
rlabel metal1 35696 55386 35696 55386 0 net9
rlabel metal2 24242 1928 24242 1928 0 net90
rlabel metal2 24518 2336 24518 2336 0 net91
rlabel metal2 24794 1418 24794 1418 0 net92
rlabel metal2 25070 1792 25070 1792 0 net93
rlabel metal2 25346 1520 25346 1520 0 net94
rlabel metal2 25622 1656 25622 1656 0 net95
rlabel metal2 25898 1622 25898 1622 0 net96
rlabel metal2 38778 2992 38778 2992 0 net97
rlabel metal2 35926 3910 35926 3910 0 net98
rlabel metal2 40066 2992 40066 2992 0 net99
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
