magic
tech sky130A
magscale 1 2
timestamp 1672273952
<< viali >>
rect 3709 57545 3743 57579
rect 5273 57545 5307 57579
rect 10793 57545 10827 57579
rect 12173 57545 12207 57579
rect 13553 57545 13587 57579
rect 14933 57545 14967 57579
rect 16313 57545 16347 57579
rect 17693 57545 17727 57579
rect 19165 57545 19199 57579
rect 20453 57545 20487 57579
rect 22109 57545 22143 57579
rect 23213 57545 23247 57579
rect 25145 57545 25179 57579
rect 26065 57545 26099 57579
rect 28089 57545 28123 57579
rect 28733 57545 28767 57579
rect 40049 57545 40083 57579
rect 4445 57477 4479 57511
rect 36093 57477 36127 57511
rect 41889 57477 41923 57511
rect 45845 57477 45879 57511
rect 52653 57477 52687 57511
rect 5457 57409 5491 57443
rect 5917 57409 5951 57443
rect 6561 57409 6595 57443
rect 7297 57409 7331 57443
rect 7941 57409 7975 57443
rect 8677 57409 8711 57443
rect 9321 57409 9355 57443
rect 10977 57409 11011 57443
rect 11437 57409 11471 57443
rect 12357 57409 12391 57443
rect 13737 57409 13771 57443
rect 14197 57409 14231 57443
rect 15117 57409 15151 57443
rect 16497 57409 16531 57443
rect 16957 57409 16991 57443
rect 17877 57409 17911 57443
rect 18337 57409 18371 57443
rect 19349 57409 19383 57443
rect 20649 57409 20683 57443
rect 22293 57409 22327 57443
rect 23397 57409 23431 57443
rect 24041 57409 24075 57443
rect 24961 57409 24995 57443
rect 25881 57409 25915 57443
rect 27169 57409 27203 57443
rect 27353 57409 27387 57443
rect 27905 57409 27939 57443
rect 28917 57409 28951 57443
rect 29469 57409 29503 57443
rect 30941 57409 30975 57443
rect 32689 57409 32723 57443
rect 33977 57409 34011 57443
rect 34161 57409 34195 57443
rect 34253 57409 34287 57443
rect 34897 57409 34931 57443
rect 35633 57409 35667 57443
rect 36737 57409 36771 57443
rect 38025 57409 38059 57443
rect 40417 57409 40451 57443
rect 42073 57409 42107 57443
rect 42901 57409 42935 57443
rect 47041 57409 47075 57443
rect 48513 57409 48547 57443
rect 49801 57409 49835 57443
rect 51457 57409 51491 57443
rect 53481 57409 53515 57443
rect 54401 57409 54435 57443
rect 55597 57409 55631 57443
rect 56057 57409 56091 57443
rect 24225 57341 24259 57375
rect 30297 57341 30331 57375
rect 32413 57341 32447 57375
rect 37013 57341 37047 57375
rect 38301 57341 38335 57375
rect 40233 57341 40267 57375
rect 40325 57341 40359 57375
rect 40509 57341 40543 57375
rect 43177 57341 43211 57375
rect 47317 57341 47351 57375
rect 48789 57341 48823 57375
rect 50077 57341 50111 57375
rect 4629 57273 4663 57307
rect 21465 57273 21499 57307
rect 29653 57273 29687 57307
rect 33793 57273 33827 57307
rect 35449 57273 35483 57307
rect 54585 57273 54619 57307
rect 23857 57205 23891 57239
rect 26709 57205 26743 57239
rect 27353 57205 27387 57239
rect 33241 57205 33275 57239
rect 34805 57205 34839 57239
rect 41061 57205 41095 57239
rect 41705 57205 41739 57239
rect 44189 57205 44223 57239
rect 44833 57205 44867 57239
rect 45753 57205 45787 57239
rect 46397 57205 46431 57239
rect 51641 57205 51675 57239
rect 52745 57205 52779 57239
rect 55413 57205 55447 57239
rect 4721 57001 4755 57035
rect 10333 57001 10367 57035
rect 13001 57001 13035 57035
rect 16313 57001 16347 57035
rect 19901 57001 19935 57035
rect 21281 57001 21315 57035
rect 23489 57001 23523 57035
rect 24593 57001 24627 57035
rect 25053 57001 25087 57035
rect 29101 57001 29135 57035
rect 30757 57001 30791 57035
rect 34253 57001 34287 57035
rect 40233 57001 40267 57035
rect 48145 57001 48179 57035
rect 49433 57001 49467 57035
rect 50721 57001 50755 57035
rect 52193 57001 52227 57035
rect 53481 57001 53515 57035
rect 54401 57001 54435 57035
rect 55045 57001 55079 57035
rect 55689 57001 55723 57035
rect 56241 57001 56275 57035
rect 11161 56933 11195 56967
rect 22937 56933 22971 56967
rect 28365 56933 28399 56967
rect 32873 56933 32907 56967
rect 33241 56933 33275 56967
rect 40601 56933 40635 56967
rect 41153 56933 41187 56967
rect 43821 56933 43855 56967
rect 47501 56933 47535 56967
rect 50077 56933 50111 56967
rect 51365 56933 51399 56967
rect 52837 56933 52871 56967
rect 27629 56865 27663 56899
rect 29561 56865 29595 56899
rect 31033 56865 31067 56899
rect 31125 56865 31159 56899
rect 35357 56865 35391 56899
rect 37749 56865 37783 56899
rect 38025 56865 38059 56899
rect 41797 56865 41831 56899
rect 42809 56865 42843 56899
rect 43729 56865 43763 56899
rect 43913 56865 43947 56899
rect 48789 56865 48823 56899
rect 23397 56797 23431 56831
rect 23916 56797 23950 56831
rect 25234 56797 25268 56831
rect 25605 56797 25639 56831
rect 25697 56797 25731 56831
rect 26433 56797 26467 56831
rect 26617 56797 26651 56831
rect 27353 56797 27387 56831
rect 27445 56797 27479 56831
rect 27721 56797 27755 56831
rect 28641 56797 28675 56831
rect 29285 56797 29319 56831
rect 29469 56797 29503 56831
rect 29653 56797 29687 56831
rect 29837 56797 29871 56831
rect 30941 56797 30975 56831
rect 31217 56797 31251 56831
rect 31922 56797 31956 56831
rect 32321 56797 32355 56831
rect 32413 56797 32447 56831
rect 33057 56797 33091 56831
rect 33333 56797 33367 56831
rect 34897 56797 34931 56831
rect 35265 56797 35299 56831
rect 36001 56797 36035 56831
rect 36277 56797 36311 56831
rect 36461 56797 36495 56831
rect 36737 56797 36771 56831
rect 37933 56797 37967 56831
rect 38117 56797 38151 56831
rect 38209 56797 38243 56831
rect 38761 56797 38795 56831
rect 40417 56797 40451 56831
rect 40693 56797 40727 56831
rect 41334 56797 41368 56831
rect 41705 56797 41739 56831
rect 42993 56797 43027 56831
rect 43177 56797 43211 56831
rect 43269 56797 43303 56831
rect 44189 56797 44223 56831
rect 44557 56797 44591 56831
rect 45201 56797 45235 56831
rect 46213 56797 46247 56831
rect 47041 56797 47075 56831
rect 27169 56729 27203 56763
rect 28365 56729 28399 56763
rect 5641 56661 5675 56695
rect 23857 56661 23891 56695
rect 24041 56661 24075 56695
rect 25237 56661 25271 56695
rect 26249 56661 26283 56695
rect 28549 56661 28583 56695
rect 31769 56661 31803 56695
rect 31953 56661 31987 56695
rect 34989 56661 35023 56695
rect 36093 56661 36127 56695
rect 38991 56661 39025 56695
rect 41337 56661 41371 56695
rect 42349 56661 42383 56695
rect 45017 56661 45051 56695
rect 46857 56661 46891 56695
rect 23489 56457 23523 56491
rect 26709 56457 26743 56491
rect 26893 56457 26927 56491
rect 27997 56457 28031 56491
rect 31493 56457 31527 56491
rect 35357 56457 35391 56491
rect 48329 56457 48363 56491
rect 49709 56457 49743 56491
rect 51273 56457 51307 56491
rect 52469 56457 52503 56491
rect 54217 56457 54251 56491
rect 35725 56389 35759 56423
rect 36645 56389 36679 56423
rect 43361 56389 43395 56423
rect 22661 56321 22695 56355
rect 23305 56321 23339 56355
rect 23949 56321 23983 56355
rect 25513 56321 25547 56355
rect 26249 56321 26283 56355
rect 26768 56321 26802 56355
rect 27353 56321 27387 56355
rect 27537 56321 27571 56355
rect 28181 56321 28215 56355
rect 28365 56321 28399 56355
rect 29101 56321 29135 56355
rect 29377 56321 29411 56355
rect 29561 56321 29595 56355
rect 30021 56321 30055 56355
rect 31677 56321 31711 56355
rect 32413 56321 32447 56355
rect 33333 56321 33367 56355
rect 33425 56321 33459 56355
rect 33609 56321 33643 56355
rect 33701 56321 33735 56355
rect 34161 56321 34195 56355
rect 34345 56321 34379 56355
rect 34621 56321 34655 56355
rect 35541 56321 35575 56355
rect 36461 56321 36495 56355
rect 36737 56321 36771 56355
rect 38761 56321 38795 56355
rect 40049 56321 40083 56355
rect 40141 56321 40175 56355
rect 40233 56321 40267 56355
rect 40371 56321 40405 56355
rect 41061 56321 41095 56355
rect 41245 56321 41279 56355
rect 41981 56321 42015 56355
rect 42165 56321 42199 56355
rect 42257 56321 42291 56355
rect 42426 56321 42460 56355
rect 42533 56321 42567 56355
rect 43269 56321 43303 56355
rect 43545 56321 43579 56355
rect 44649 56321 44683 56355
rect 45568 56321 45602 56355
rect 45661 56321 45695 56355
rect 47409 56321 47443 56355
rect 24225 56253 24259 56287
rect 25329 56253 25363 56287
rect 28917 56253 28951 56287
rect 29285 56253 29319 56287
rect 31953 56253 31987 56287
rect 38117 56253 38151 56287
rect 38577 56253 38611 56287
rect 38945 56253 38979 56287
rect 40509 56253 40543 56287
rect 41521 56253 41555 56287
rect 44557 56253 44591 56287
rect 46765 56253 46799 56287
rect 26341 56185 26375 56219
rect 27537 56185 27571 56219
rect 29193 56185 29227 56219
rect 36277 56185 36311 56219
rect 37841 56185 37875 56219
rect 43729 56185 43763 56219
rect 46121 56185 46155 56219
rect 22109 56117 22143 56151
rect 25697 56117 25731 56151
rect 30665 56117 30699 56151
rect 31861 56117 31895 56151
rect 33149 56117 33183 56151
rect 34529 56117 34563 56151
rect 37657 56117 37691 56151
rect 39865 56117 39899 56151
rect 41429 56117 41463 56151
rect 44373 56117 44407 56151
rect 45477 56117 45511 56151
rect 24777 55913 24811 55947
rect 26249 55913 26283 55947
rect 27721 55913 27755 55947
rect 35725 55913 35759 55947
rect 36829 55913 36863 55947
rect 38117 55913 38151 55947
rect 40233 55913 40267 55947
rect 41429 55913 41463 55947
rect 42349 55913 42383 55947
rect 42717 55913 42751 55947
rect 44649 55913 44683 55947
rect 46765 55913 46799 55947
rect 47317 55913 47351 55947
rect 31493 55845 31527 55879
rect 34713 55845 34747 55879
rect 37381 55845 37415 55879
rect 44189 55845 44223 55879
rect 45017 55845 45051 55879
rect 46305 55845 46339 55879
rect 23213 55777 23247 55811
rect 23673 55777 23707 55811
rect 28457 55777 28491 55811
rect 28733 55777 28767 55811
rect 28917 55777 28951 55811
rect 34989 55777 35023 55811
rect 36645 55777 36679 55811
rect 43269 55777 43303 55811
rect 23857 55709 23891 55743
rect 24593 55709 24627 55743
rect 25237 55709 25271 55743
rect 25421 55709 25455 55743
rect 25605 55709 25639 55743
rect 26065 55709 26099 55743
rect 26709 55709 26743 55743
rect 26893 55709 26927 55743
rect 26985 55709 27019 55743
rect 27537 55709 27571 55743
rect 28641 55709 28675 55743
rect 28825 55709 28859 55743
rect 29653 55709 29687 55743
rect 29837 55709 29871 55743
rect 30849 55709 30883 55743
rect 31309 55709 31343 55743
rect 32137 55709 32171 55743
rect 32413 55709 32447 55743
rect 33057 55709 33091 55743
rect 33241 55709 33275 55743
rect 33333 55709 33367 55743
rect 35081 55709 35115 55743
rect 36553 55709 36587 55743
rect 37565 55709 37599 55743
rect 37657 55709 37691 55743
rect 38301 55709 38335 55743
rect 38393 55709 38427 55743
rect 38577 55709 38611 55743
rect 38669 55709 38703 55743
rect 39313 55709 39347 55743
rect 39497 55709 39531 55743
rect 41061 55709 41095 55743
rect 42533 55709 42567 55743
rect 42809 55709 42843 55743
rect 43913 55709 43947 55743
rect 44005 55709 44039 55743
rect 44189 55709 44223 55743
rect 44833 55709 44867 55743
rect 44925 55709 44959 55743
rect 45109 55709 45143 55743
rect 30987 55641 31021 55675
rect 31125 55641 31159 55675
rect 31217 55641 31251 55675
rect 31953 55641 31987 55675
rect 32873 55641 32907 55675
rect 37381 55641 37415 55675
rect 39129 55641 39163 55675
rect 40417 55641 40451 55675
rect 40601 55641 40635 55675
rect 41245 55641 41279 55675
rect 24041 55573 24075 55607
rect 29469 55573 29503 55607
rect 30389 55573 30423 55607
rect 32321 55573 32355 55607
rect 23857 55369 23891 55403
rect 25513 55369 25547 55403
rect 26249 55369 26283 55403
rect 30757 55369 30791 55403
rect 33057 55369 33091 55403
rect 34430 55369 34464 55403
rect 34989 55369 35023 55403
rect 38117 55369 38151 55403
rect 38485 55369 38519 55403
rect 40042 55369 40076 55403
rect 44465 55369 44499 55403
rect 45109 55369 45143 55403
rect 45569 55369 45603 55403
rect 29009 55301 29043 55335
rect 29745 55301 29779 55335
rect 29929 55301 29963 55335
rect 33609 55301 33643 55335
rect 34345 55301 34379 55335
rect 34529 55301 34563 55335
rect 39037 55301 39071 55335
rect 39957 55301 39991 55335
rect 40141 55301 40175 55335
rect 44005 55301 44039 55335
rect 24041 55233 24075 55267
rect 25697 55233 25731 55267
rect 26433 55233 26467 55267
rect 26893 55233 26927 55267
rect 26985 55233 27019 55267
rect 27537 55233 27571 55267
rect 27721 55233 27755 55267
rect 27813 55233 27847 55267
rect 29561 55233 29595 55267
rect 30389 55233 30423 55267
rect 30573 55233 30607 55267
rect 31769 55233 31803 55267
rect 32689 55233 32723 55267
rect 32873 55233 32907 55267
rect 33701 55233 33735 55267
rect 34253 55233 34287 55267
rect 35173 55233 35207 55267
rect 35357 55233 35391 55267
rect 35449 55233 35483 55267
rect 36276 55233 36310 55267
rect 36369 55233 36403 55267
rect 38301 55233 38335 55267
rect 38577 55233 38611 55267
rect 39221 55233 39255 55267
rect 39865 55233 39899 55267
rect 40693 55233 40727 55267
rect 42073 55233 42107 55267
rect 36001 55165 36035 55199
rect 37289 55165 37323 55199
rect 39405 55165 39439 55199
rect 42533 55165 42567 55199
rect 43269 55165 43303 55199
rect 28641 55097 28675 55131
rect 35265 55097 35299 55131
rect 24777 55029 24811 55063
rect 27629 55029 27663 55063
rect 28549 55029 28583 55063
rect 31861 55029 31895 55063
rect 32229 55029 32263 55063
rect 40785 55029 40819 55063
rect 41153 55029 41187 55063
rect 41613 55029 41647 55063
rect 41889 55029 41923 55063
rect 25789 54825 25823 54859
rect 26249 54825 26283 54859
rect 26801 54825 26835 54859
rect 27721 54825 27755 54859
rect 29101 54825 29135 54859
rect 30113 54825 30147 54859
rect 31033 54825 31067 54859
rect 35173 54825 35207 54859
rect 35817 54825 35851 54859
rect 36461 54825 36495 54859
rect 37197 54825 37231 54859
rect 37841 54825 37875 54859
rect 38485 54825 38519 54859
rect 39589 54825 39623 54859
rect 41705 54825 41739 54859
rect 44925 54825 44959 54859
rect 24409 54757 24443 54791
rect 25237 54757 25271 54791
rect 28641 54757 28675 54791
rect 43545 54757 43579 54791
rect 39313 54689 39347 54723
rect 40785 54689 40819 54723
rect 44005 54689 44039 54723
rect 44557 54689 44591 54723
rect 45017 54689 45051 54723
rect 28365 54621 28399 54655
rect 29277 54631 29311 54665
rect 29369 54621 29403 54655
rect 29546 54621 29580 54655
rect 29653 54621 29687 54655
rect 30757 54621 30791 54655
rect 31953 54621 31987 54655
rect 32137 54621 32171 54655
rect 32413 54621 32447 54655
rect 33057 54621 33091 54655
rect 33333 54621 33367 54655
rect 34437 54621 34471 54655
rect 34529 54621 34563 54655
rect 34621 54621 34655 54655
rect 39221 54621 39255 54655
rect 40969 54621 41003 54655
rect 41245 54621 41279 54655
rect 42625 54621 42659 54655
rect 42717 54621 42751 54655
rect 43913 54621 43947 54655
rect 44741 54621 44775 54655
rect 28641 54553 28675 54587
rect 30849 54553 30883 54587
rect 31033 54553 31067 54587
rect 40233 54553 40267 54587
rect 41153 54553 41187 54587
rect 28457 54485 28491 54519
rect 32321 54485 32355 54519
rect 32873 54485 32907 54519
rect 33241 54485 33275 54519
rect 34253 54485 34287 54519
rect 42441 54485 42475 54519
rect 43085 54485 43119 54519
rect 27261 54281 27295 54315
rect 27905 54281 27939 54315
rect 28917 54281 28951 54315
rect 29377 54281 29411 54315
rect 32781 54281 32815 54315
rect 33609 54281 33643 54315
rect 34253 54281 34287 54315
rect 36645 54281 36679 54315
rect 37289 54281 37323 54315
rect 39037 54281 39071 54315
rect 40325 54281 40359 54315
rect 41521 54281 41555 54315
rect 41981 54281 42015 54315
rect 39681 54213 39715 54247
rect 42349 54213 42383 54247
rect 43269 54213 43303 54247
rect 28549 54145 28583 54179
rect 29561 54145 29595 54179
rect 30389 54145 30423 54179
rect 32413 54145 32447 54179
rect 33793 54145 33827 54179
rect 35003 54145 35037 54179
rect 35725 54145 35759 54179
rect 36001 54145 36035 54179
rect 38301 54145 38335 54179
rect 39129 54145 39163 54179
rect 40141 54145 40175 54179
rect 41153 54145 41187 54179
rect 42165 54145 42199 54179
rect 42441 54145 42475 54179
rect 43453 54145 43487 54179
rect 43545 54145 43579 54179
rect 43637 54145 43671 54179
rect 28457 54077 28491 54111
rect 29745 54077 29779 54111
rect 30481 54077 30515 54111
rect 30757 54077 30791 54111
rect 32321 54077 32355 54111
rect 33885 54077 33919 54111
rect 35173 54077 35207 54111
rect 41245 54077 41279 54111
rect 26617 54009 26651 54043
rect 34713 54009 34747 54043
rect 36185 54009 36219 54043
rect 31401 53941 31435 53975
rect 35817 53941 35851 53975
rect 29837 53737 29871 53771
rect 32413 53737 32447 53771
rect 32597 53737 32631 53771
rect 33333 53737 33367 53771
rect 33517 53737 33551 53771
rect 34897 53737 34931 53771
rect 35449 53737 35483 53771
rect 35909 53737 35943 53771
rect 40233 53737 40267 53771
rect 41889 53737 41923 53771
rect 42073 53737 42107 53771
rect 27537 53669 27571 53703
rect 29193 53669 29227 53703
rect 34345 53669 34379 53703
rect 40785 53601 40819 53635
rect 41337 53601 41371 53635
rect 30021 53533 30055 53567
rect 30205 53533 30239 53567
rect 32873 53533 32907 53567
rect 33485 53465 33519 53499
rect 33701 53465 33735 53499
rect 42257 53465 42291 53499
rect 28641 53397 28675 53431
rect 42057 53397 42091 53431
rect 33701 53193 33735 53227
rect 35357 53193 35391 53227
rect 40785 53193 40819 53227
rect 32597 53125 32631 53159
rect 33241 53125 33275 53159
rect 34345 53125 34379 53159
rect 34897 53125 34931 53159
rect 34253 52037 34287 52071
rect 34069 51901 34103 51935
rect 35817 51901 35851 51935
rect 34253 51561 34287 51595
rect 30021 8449 30055 8483
rect 30113 8313 30147 8347
rect 29009 8041 29043 8075
rect 29469 7837 29503 7871
rect 30113 7837 30147 7871
rect 30849 7837 30883 7871
rect 30941 7701 30975 7735
rect 26985 7361 27019 7395
rect 30021 7361 30055 7395
rect 32137 7361 32171 7395
rect 27721 7293 27755 7327
rect 27905 7293 27939 7327
rect 29193 7293 29227 7327
rect 30205 7293 30239 7327
rect 26893 7157 26927 7191
rect 31309 7157 31343 7191
rect 32229 7157 32263 7191
rect 28733 6817 28767 6851
rect 30297 6817 30331 6851
rect 31217 6817 31251 6851
rect 31493 6817 31527 6851
rect 26893 6749 26927 6783
rect 27721 6749 27755 6783
rect 31033 6749 31067 6783
rect 34253 6749 34287 6783
rect 28917 6681 28951 6715
rect 26433 6613 26467 6647
rect 26985 6613 27019 6647
rect 34345 6613 34379 6647
rect 27813 6341 27847 6375
rect 30573 6341 30607 6375
rect 26709 6273 26743 6307
rect 27629 6273 27663 6307
rect 30297 6273 30331 6307
rect 31309 6273 31343 6307
rect 26985 6205 27019 6239
rect 28089 6205 28123 6239
rect 32597 6205 32631 6239
rect 33517 6205 33551 6239
rect 33701 6205 33735 6239
rect 26249 6137 26283 6171
rect 25329 6069 25363 6103
rect 34345 6069 34379 6103
rect 29469 5865 29503 5899
rect 32505 5865 32539 5899
rect 33057 5865 33091 5899
rect 26065 5729 26099 5763
rect 27537 5729 27571 5763
rect 30021 5729 30055 5763
rect 30205 5729 30239 5763
rect 30573 5729 30607 5763
rect 34253 5729 34287 5763
rect 34437 5729 34471 5763
rect 34713 5729 34747 5763
rect 24133 5661 24167 5695
rect 24593 5661 24627 5695
rect 25421 5661 25455 5695
rect 25881 5661 25915 5695
rect 28917 5661 28951 5695
rect 29561 5661 29595 5695
rect 32965 5661 32999 5695
rect 24685 5525 24719 5559
rect 27721 5321 27755 5355
rect 25513 5253 25547 5287
rect 31493 5253 31527 5287
rect 33793 5253 33827 5287
rect 25329 5185 25363 5219
rect 27629 5185 27663 5219
rect 28273 5185 28307 5219
rect 28917 5185 28951 5219
rect 24133 5117 24167 5151
rect 26249 5117 26283 5151
rect 28365 5117 28399 5151
rect 29101 5117 29135 5151
rect 30389 5117 30423 5151
rect 31309 5117 31343 5151
rect 31769 5117 31803 5151
rect 33609 5117 33643 5151
rect 34069 5117 34103 5151
rect 23213 4981 23247 5015
rect 24777 4981 24811 5015
rect 36093 4981 36127 5015
rect 24777 4777 24811 4811
rect 32781 4777 32815 4811
rect 23489 4709 23523 4743
rect 25421 4709 25455 4743
rect 25881 4641 25915 4675
rect 26433 4641 26467 4675
rect 30757 4641 30791 4675
rect 36093 4641 36127 4675
rect 21557 4573 21591 4607
rect 22661 4573 22695 4607
rect 23949 4573 23983 4607
rect 28549 4573 28583 4607
rect 29009 4573 29043 4607
rect 29837 4573 29871 4607
rect 30297 4573 30331 4607
rect 33425 4573 33459 4607
rect 36737 4573 36771 4607
rect 24041 4505 24075 4539
rect 26065 4505 26099 4539
rect 29101 4505 29135 4539
rect 30481 4505 30515 4539
rect 34253 4505 34287 4539
rect 35909 4505 35943 4539
rect 36645 4505 36679 4539
rect 34345 4165 34379 4199
rect 23949 4097 23983 4131
rect 24593 4097 24627 4131
rect 25329 4097 25363 4131
rect 25973 4097 26007 4131
rect 28917 4097 28951 4131
rect 31309 4097 31343 4131
rect 34529 4097 34563 4131
rect 35081 4097 35115 4131
rect 35173 4097 35207 4131
rect 23489 4029 23523 4063
rect 26617 4029 26651 4063
rect 26801 4029 26835 4063
rect 28457 4029 28491 4063
rect 29101 4029 29135 4063
rect 29745 4029 29779 4063
rect 33057 4029 33091 4063
rect 22201 3961 22235 3995
rect 24041 3961 24075 3995
rect 37933 3961 37967 3995
rect 19901 3893 19935 3927
rect 20729 3893 20763 3927
rect 21557 3893 21591 3927
rect 22845 3893 22879 3927
rect 24685 3893 24719 3927
rect 25421 3893 25455 3927
rect 26065 3893 26099 3927
rect 31953 3893 31987 3927
rect 35633 3893 35667 3927
rect 36277 3893 36311 3927
rect 37289 3893 37323 3927
rect 38669 3893 38703 3927
rect 30849 3689 30883 3723
rect 37841 3689 37875 3723
rect 21097 3621 21131 3655
rect 37197 3621 37231 3655
rect 40877 3621 40911 3655
rect 23029 3553 23063 3587
rect 26065 3553 26099 3587
rect 28457 3553 28491 3587
rect 28733 3553 28767 3587
rect 31493 3553 31527 3587
rect 31953 3553 31987 3587
rect 34437 3553 34471 3587
rect 36093 3553 36127 3587
rect 39129 3553 39163 3587
rect 41521 3553 41555 3587
rect 9413 3485 9447 3519
rect 10885 3485 10919 3519
rect 12541 3485 12575 3519
rect 13645 3485 13679 3519
rect 14749 3485 14783 3519
rect 15577 3485 15611 3519
rect 16681 3485 16715 3519
rect 17417 3485 17451 3519
rect 18245 3485 18279 3519
rect 18981 3485 19015 3519
rect 19809 3485 19843 3519
rect 20453 3485 20487 3519
rect 21741 3485 21775 3519
rect 22293 3485 22327 3519
rect 22937 3485 22971 3519
rect 23581 3485 23615 3519
rect 25881 3485 25915 3519
rect 28273 3485 28307 3519
rect 30757 3485 30791 3519
rect 36737 3485 36771 3519
rect 38485 3485 38519 3519
rect 40233 3485 40267 3519
rect 42165 3485 42199 3519
rect 42809 3485 42843 3519
rect 43453 3485 43487 3519
rect 44189 3485 44223 3519
rect 46213 3485 46247 3519
rect 46857 3485 46891 3519
rect 48329 3485 48363 3519
rect 49433 3485 49467 3519
rect 50261 3485 50295 3519
rect 52193 3485 52227 3519
rect 22385 3417 22419 3451
rect 23765 3417 23799 3451
rect 25421 3417 25455 3451
rect 27721 3417 27755 3451
rect 31677 3417 31711 3451
rect 35909 3417 35943 3451
rect 36645 3349 36679 3383
rect 30665 3145 30699 3179
rect 23397 3077 23431 3111
rect 25789 3077 25823 3111
rect 28089 3077 28123 3111
rect 33241 3077 33275 3111
rect 35541 3077 35575 3111
rect 37381 3077 37415 3111
rect 20913 3009 20947 3043
rect 22201 3009 22235 3043
rect 22845 3009 22879 3043
rect 23489 3009 23523 3043
rect 24593 3009 24627 3043
rect 27905 3009 27939 3043
rect 30573 3009 30607 3043
rect 33425 3009 33459 3043
rect 35725 3009 35759 3043
rect 37289 3009 37323 3043
rect 39865 3009 39899 3043
rect 41797 3009 41831 3043
rect 16221 2941 16255 2975
rect 19625 2941 19659 2975
rect 24685 2941 24719 2975
rect 25605 2941 25639 2975
rect 27445 2941 27479 2975
rect 28641 2941 28675 2975
rect 32229 2941 32263 2975
rect 33885 2941 33919 2975
rect 37933 2941 37967 2975
rect 41153 2941 41187 2975
rect 46489 2941 46523 2975
rect 47777 2941 47811 2975
rect 20269 2873 20303 2907
rect 22109 2873 22143 2907
rect 24133 2873 24167 2907
rect 38577 2873 38611 2907
rect 40509 2873 40543 2907
rect 42441 2873 42475 2907
rect 43913 2873 43947 2907
rect 45201 2873 45235 2907
rect 48421 2873 48455 2907
rect 49893 2873 49927 2907
rect 51825 2873 51859 2907
rect 53113 2873 53147 2907
rect 7757 2805 7791 2839
rect 8677 2805 8711 2839
rect 9597 2805 9631 2839
rect 10241 2805 10275 2839
rect 10885 2805 10919 2839
rect 11529 2805 11563 2839
rect 12173 2805 12207 2839
rect 12817 2805 12851 2839
rect 13645 2805 13679 2839
rect 14289 2805 14323 2839
rect 14933 2805 14967 2839
rect 15577 2805 15611 2839
rect 16865 2805 16899 2839
rect 17509 2805 17543 2839
rect 18153 2805 18187 2839
rect 18797 2805 18831 2839
rect 21557 2805 21591 2839
rect 36185 2805 36219 2839
rect 39221 2805 39255 2839
rect 43269 2805 43303 2839
rect 44557 2805 44591 2839
rect 45845 2805 45879 2839
rect 47133 2805 47167 2839
rect 49249 2805 49283 2839
rect 50537 2805 50571 2839
rect 51181 2805 51215 2839
rect 52469 2805 52503 2839
rect 22477 2601 22511 2635
rect 23765 2601 23799 2635
rect 37473 2601 37507 2635
rect 38669 2601 38703 2635
rect 49801 2601 49835 2635
rect 9045 2533 9079 2567
rect 10701 2533 10735 2567
rect 14289 2533 14323 2567
rect 17233 2533 17267 2567
rect 18521 2533 18555 2567
rect 20821 2533 20855 2567
rect 38025 2533 38059 2567
rect 40969 2533 41003 2567
rect 43269 2533 43303 2567
rect 46857 2533 46891 2567
rect 50445 2533 50479 2567
rect 52101 2533 52135 2567
rect 11989 2465 12023 2499
rect 16589 2465 16623 2499
rect 17877 2465 17911 2499
rect 19533 2465 19567 2499
rect 23121 2465 23155 2499
rect 25513 2465 25547 2499
rect 28457 2465 28491 2499
rect 29469 2465 29503 2499
rect 31125 2465 31159 2499
rect 32505 2465 32539 2499
rect 32689 2465 32723 2499
rect 43913 2465 43947 2499
rect 46213 2465 46247 2499
rect 48513 2465 48547 2499
rect 51457 2465 51491 2499
rect 53389 2465 53423 2499
rect 7757 2397 7791 2431
rect 8401 2397 8435 2431
rect 9689 2397 9723 2431
rect 11345 2397 11379 2431
rect 12633 2397 12667 2431
rect 13645 2397 13679 2431
rect 14933 2397 14967 2431
rect 15577 2397 15611 2431
rect 20177 2397 20211 2431
rect 21465 2397 21499 2431
rect 24225 2397 24259 2431
rect 35633 2397 35667 2431
rect 36921 2397 36955 2431
rect 37381 2397 37415 2431
rect 39681 2397 39715 2431
rect 40325 2397 40359 2431
rect 41613 2397 41647 2431
rect 42625 2397 42659 2431
rect 44557 2397 44591 2431
rect 45569 2397 45603 2431
rect 47501 2397 47535 2431
rect 49157 2397 49191 2431
rect 52745 2397 52779 2431
rect 25697 2329 25731 2363
rect 27353 2329 27387 2363
rect 28641 2329 28675 2363
rect 33793 2329 33827 2363
rect 35449 2329 35483 2363
rect 36829 2329 36863 2363
rect 24317 2261 24351 2295
<< metal1 >>
rect 23198 57944 23204 57996
rect 23256 57984 23262 57996
rect 23256 57956 25176 57984
rect 23256 57944 23262 57956
rect 15102 57876 15108 57928
rect 15160 57916 15166 57928
rect 25038 57916 25044 57928
rect 15160 57888 25044 57916
rect 15160 57876 15166 57888
rect 25038 57876 25044 57888
rect 25096 57876 25102 57928
rect 25148 57916 25176 57956
rect 25148 57888 27108 57916
rect 27080 57860 27108 57888
rect 12342 57808 12348 57860
rect 12400 57848 12406 57860
rect 26970 57848 26976 57860
rect 12400 57820 26976 57848
rect 12400 57808 12406 57820
rect 26970 57808 26976 57820
rect 27028 57808 27034 57860
rect 27062 57808 27068 57860
rect 27120 57848 27126 57860
rect 33686 57848 33692 57860
rect 27120 57820 33692 57848
rect 27120 57808 27126 57820
rect 33686 57808 33692 57820
rect 33744 57808 33750 57860
rect 23750 57740 23756 57792
rect 23808 57780 23814 57792
rect 39942 57780 39948 57792
rect 23808 57752 39948 57780
rect 23808 57740 23814 57752
rect 39942 57740 39948 57752
rect 40000 57740 40006 57792
rect 41414 57740 41420 57792
rect 41472 57780 41478 57792
rect 45186 57780 45192 57792
rect 41472 57752 45192 57780
rect 41472 57740 41478 57752
rect 45186 57740 45192 57752
rect 45244 57740 45250 57792
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 3694 57576 3700 57588
rect 3655 57548 3700 57576
rect 3694 57536 3700 57548
rect 3752 57576 3758 57588
rect 3752 57548 4476 57576
rect 3752 57536 3758 57548
rect 4448 57517 4476 57548
rect 5074 57536 5080 57588
rect 5132 57576 5138 57588
rect 5261 57579 5319 57585
rect 5261 57576 5273 57579
rect 5132 57548 5273 57576
rect 5132 57536 5138 57548
rect 5261 57545 5273 57548
rect 5307 57545 5319 57579
rect 5261 57539 5319 57545
rect 10594 57536 10600 57588
rect 10652 57576 10658 57588
rect 10781 57579 10839 57585
rect 10781 57576 10793 57579
rect 10652 57548 10793 57576
rect 10652 57536 10658 57548
rect 10781 57545 10793 57548
rect 10827 57545 10839 57579
rect 10781 57539 10839 57545
rect 11974 57536 11980 57588
rect 12032 57576 12038 57588
rect 12161 57579 12219 57585
rect 12161 57576 12173 57579
rect 12032 57548 12173 57576
rect 12032 57536 12038 57548
rect 12161 57545 12173 57548
rect 12207 57545 12219 57579
rect 12161 57539 12219 57545
rect 13354 57536 13360 57588
rect 13412 57576 13418 57588
rect 13541 57579 13599 57585
rect 13541 57576 13553 57579
rect 13412 57548 13553 57576
rect 13412 57536 13418 57548
rect 13541 57545 13553 57548
rect 13587 57545 13599 57579
rect 13541 57539 13599 57545
rect 14734 57536 14740 57588
rect 14792 57576 14798 57588
rect 14921 57579 14979 57585
rect 14921 57576 14933 57579
rect 14792 57548 14933 57576
rect 14792 57536 14798 57548
rect 14921 57545 14933 57548
rect 14967 57545 14979 57579
rect 14921 57539 14979 57545
rect 16114 57536 16120 57588
rect 16172 57576 16178 57588
rect 16301 57579 16359 57585
rect 16301 57576 16313 57579
rect 16172 57548 16313 57576
rect 16172 57536 16178 57548
rect 16301 57545 16313 57548
rect 16347 57545 16359 57579
rect 16301 57539 16359 57545
rect 17494 57536 17500 57588
rect 17552 57576 17558 57588
rect 17681 57579 17739 57585
rect 17681 57576 17693 57579
rect 17552 57548 17693 57576
rect 17552 57536 17558 57548
rect 17681 57545 17693 57548
rect 17727 57545 17739 57579
rect 17681 57539 17739 57545
rect 18874 57536 18880 57588
rect 18932 57576 18938 57588
rect 19153 57579 19211 57585
rect 19153 57576 19165 57579
rect 18932 57548 19165 57576
rect 18932 57536 18938 57548
rect 19153 57545 19165 57548
rect 19199 57545 19211 57579
rect 19153 57539 19211 57545
rect 20254 57536 20260 57588
rect 20312 57576 20318 57588
rect 20441 57579 20499 57585
rect 20441 57576 20453 57579
rect 20312 57548 20453 57576
rect 20312 57536 20318 57548
rect 20441 57545 20453 57548
rect 20487 57545 20499 57579
rect 20441 57539 20499 57545
rect 22094 57536 22100 57588
rect 22152 57576 22158 57588
rect 22152 57548 22197 57576
rect 22152 57536 22158 57548
rect 23014 57536 23020 57588
rect 23072 57576 23078 57588
rect 23201 57579 23259 57585
rect 23201 57576 23213 57579
rect 23072 57548 23213 57576
rect 23072 57536 23078 57548
rect 23201 57545 23213 57548
rect 23247 57545 23259 57579
rect 23201 57539 23259 57545
rect 24854 57536 24860 57588
rect 24912 57576 24918 57588
rect 25133 57579 25191 57585
rect 25133 57576 25145 57579
rect 24912 57548 25145 57576
rect 24912 57536 24918 57548
rect 25133 57545 25145 57548
rect 25179 57545 25191 57579
rect 25133 57539 25191 57545
rect 25774 57536 25780 57588
rect 25832 57576 25838 57588
rect 26053 57579 26111 57585
rect 26053 57576 26065 57579
rect 25832 57548 26065 57576
rect 25832 57536 25838 57548
rect 26053 57545 26065 57548
rect 26099 57545 26111 57579
rect 26053 57539 26111 57545
rect 27154 57536 27160 57588
rect 27212 57576 27218 57588
rect 28077 57579 28135 57585
rect 28077 57576 28089 57579
rect 27212 57548 28089 57576
rect 27212 57536 27218 57548
rect 28077 57545 28089 57548
rect 28123 57545 28135 57579
rect 28077 57539 28135 57545
rect 28534 57536 28540 57588
rect 28592 57576 28598 57588
rect 28721 57579 28779 57585
rect 28721 57576 28733 57579
rect 28592 57548 28733 57576
rect 28592 57536 28598 57548
rect 28721 57545 28733 57548
rect 28767 57545 28779 57579
rect 28721 57539 28779 57545
rect 33134 57536 33140 57588
rect 33192 57576 33198 57588
rect 35618 57576 35624 57588
rect 33192 57548 35624 57576
rect 33192 57536 33198 57548
rect 35618 57536 35624 57548
rect 35676 57536 35682 57588
rect 39942 57536 39948 57588
rect 40000 57576 40006 57588
rect 40037 57579 40095 57585
rect 40037 57576 40049 57579
rect 40000 57548 40049 57576
rect 40000 57536 40006 57548
rect 40037 57545 40049 57548
rect 40083 57545 40095 57579
rect 42150 57576 42156 57588
rect 40037 57539 40095 57545
rect 41892 57548 42156 57576
rect 4433 57511 4491 57517
rect 4433 57477 4445 57511
rect 4479 57477 4491 57511
rect 4433 57471 4491 57477
rect 13740 57480 21404 57508
rect 5442 57440 5448 57452
rect 5403 57412 5448 57440
rect 5442 57400 5448 57412
rect 5500 57400 5506 57452
rect 5905 57443 5963 57449
rect 5905 57409 5917 57443
rect 5951 57440 5963 57443
rect 5994 57440 6000 57452
rect 5951 57412 6000 57440
rect 5951 57409 5963 57412
rect 5905 57403 5963 57409
rect 5994 57400 6000 57412
rect 6052 57400 6058 57452
rect 6454 57400 6460 57452
rect 6512 57440 6518 57452
rect 6549 57443 6607 57449
rect 6549 57440 6561 57443
rect 6512 57412 6561 57440
rect 6512 57400 6518 57412
rect 6549 57409 6561 57412
rect 6595 57409 6607 57443
rect 6549 57403 6607 57409
rect 7285 57443 7343 57449
rect 7285 57409 7297 57443
rect 7331 57440 7343 57443
rect 7374 57440 7380 57452
rect 7331 57412 7380 57440
rect 7331 57409 7343 57412
rect 7285 57403 7343 57409
rect 7374 57400 7380 57412
rect 7432 57400 7438 57452
rect 7834 57400 7840 57452
rect 7892 57440 7898 57452
rect 7929 57443 7987 57449
rect 7929 57440 7941 57443
rect 7892 57412 7941 57440
rect 7892 57400 7898 57412
rect 7929 57409 7941 57412
rect 7975 57409 7987 57443
rect 7929 57403 7987 57409
rect 8665 57443 8723 57449
rect 8665 57409 8677 57443
rect 8711 57440 8723 57443
rect 8754 57440 8760 57452
rect 8711 57412 8760 57440
rect 8711 57409 8723 57412
rect 8665 57403 8723 57409
rect 8754 57400 8760 57412
rect 8812 57400 8818 57452
rect 9214 57400 9220 57452
rect 9272 57440 9278 57452
rect 9309 57443 9367 57449
rect 9309 57440 9321 57443
rect 9272 57412 9321 57440
rect 9272 57400 9278 57412
rect 9309 57409 9321 57412
rect 9355 57409 9367 57443
rect 10962 57440 10968 57452
rect 10923 57412 10968 57440
rect 9309 57403 9367 57409
rect 10962 57400 10968 57412
rect 11020 57400 11026 57452
rect 11425 57443 11483 57449
rect 11425 57409 11437 57443
rect 11471 57440 11483 57443
rect 11514 57440 11520 57452
rect 11471 57412 11520 57440
rect 11471 57409 11483 57412
rect 11425 57403 11483 57409
rect 11514 57400 11520 57412
rect 11572 57400 11578 57452
rect 12342 57440 12348 57452
rect 12303 57412 12348 57440
rect 12342 57400 12348 57412
rect 12400 57400 12406 57452
rect 13740 57449 13768 57480
rect 13725 57443 13783 57449
rect 13725 57409 13737 57443
rect 13771 57409 13783 57443
rect 13725 57403 13783 57409
rect 14185 57443 14243 57449
rect 14185 57409 14197 57443
rect 14231 57440 14243 57443
rect 14274 57440 14280 57452
rect 14231 57412 14280 57440
rect 14231 57409 14243 57412
rect 14185 57403 14243 57409
rect 14274 57400 14280 57412
rect 14332 57400 14338 57452
rect 15102 57440 15108 57452
rect 15063 57412 15108 57440
rect 15102 57400 15108 57412
rect 15160 57400 15166 57452
rect 16482 57440 16488 57452
rect 16443 57412 16488 57440
rect 16482 57400 16488 57412
rect 16540 57400 16546 57452
rect 16945 57443 17003 57449
rect 16945 57409 16957 57443
rect 16991 57440 17003 57443
rect 17034 57440 17040 57452
rect 16991 57412 17040 57440
rect 16991 57409 17003 57412
rect 16945 57403 17003 57409
rect 17034 57400 17040 57412
rect 17092 57400 17098 57452
rect 17862 57440 17868 57452
rect 17823 57412 17868 57440
rect 17862 57400 17868 57412
rect 17920 57400 17926 57452
rect 18325 57443 18383 57449
rect 18325 57409 18337 57443
rect 18371 57440 18383 57443
rect 18414 57440 18420 57452
rect 18371 57412 18420 57440
rect 18371 57409 18383 57412
rect 18325 57403 18383 57409
rect 18414 57400 18420 57412
rect 18472 57400 18478 57452
rect 19337 57443 19395 57449
rect 19337 57409 19349 57443
rect 19383 57440 19395 57443
rect 19383 57412 20576 57440
rect 19383 57409 19395 57412
rect 19337 57403 19395 57409
rect 4617 57307 4675 57313
rect 4617 57273 4629 57307
rect 4663 57304 4675 57307
rect 5350 57304 5356 57316
rect 4663 57276 5356 57304
rect 4663 57273 4675 57276
rect 4617 57267 4675 57273
rect 5350 57264 5356 57276
rect 5408 57264 5414 57316
rect 20548 57304 20576 57412
rect 20622 57400 20628 57452
rect 20680 57449 20686 57452
rect 20680 57443 20695 57449
rect 20683 57409 20695 57443
rect 21376 57440 21404 57480
rect 27080 57480 29500 57508
rect 21376 57412 22232 57440
rect 20680 57403 20695 57409
rect 20680 57400 20686 57403
rect 22204 57372 22232 57412
rect 22278 57400 22284 57452
rect 22336 57440 22342 57452
rect 22336 57412 22381 57440
rect 22336 57400 22342 57412
rect 23382 57400 23388 57452
rect 23440 57440 23446 57452
rect 24026 57440 24032 57452
rect 23440 57412 23485 57440
rect 23939 57412 24032 57440
rect 23440 57400 23446 57412
rect 24026 57400 24032 57412
rect 24084 57400 24090 57452
rect 24118 57400 24124 57452
rect 24176 57440 24182 57452
rect 24949 57443 25007 57449
rect 24949 57440 24961 57443
rect 24176 57412 24961 57440
rect 24176 57400 24182 57412
rect 24949 57409 24961 57412
rect 24995 57409 25007 57443
rect 24949 57403 25007 57409
rect 25590 57400 25596 57452
rect 25648 57440 25654 57452
rect 25869 57443 25927 57449
rect 25869 57440 25881 57443
rect 25648 57412 25881 57440
rect 25648 57400 25654 57412
rect 25869 57409 25881 57412
rect 25915 57409 25927 57443
rect 27080 57440 27108 57480
rect 25869 57403 25927 57409
rect 26252 57412 27108 57440
rect 23934 57372 23940 57384
rect 20824 57344 22094 57372
rect 22204 57344 23940 57372
rect 20824 57304 20852 57344
rect 21450 57304 21456 57316
rect 20548 57276 20852 57304
rect 21411 57276 21456 57304
rect 21450 57264 21456 57276
rect 21508 57264 21514 57316
rect 22066 57304 22094 57344
rect 23934 57332 23940 57344
rect 23992 57332 23998 57384
rect 23382 57304 23388 57316
rect 22066 57276 23388 57304
rect 23382 57264 23388 57276
rect 23440 57264 23446 57316
rect 24044 57304 24072 57400
rect 24213 57375 24271 57381
rect 24213 57341 24225 57375
rect 24259 57372 24271 57375
rect 24302 57372 24308 57384
rect 24259 57344 24308 57372
rect 24259 57341 24271 57344
rect 24213 57335 24271 57341
rect 24302 57332 24308 57344
rect 24360 57332 24366 57384
rect 24578 57332 24584 57384
rect 24636 57372 24642 57384
rect 26252 57372 26280 57412
rect 27154 57400 27160 57452
rect 27212 57440 27218 57452
rect 27341 57443 27399 57449
rect 27212 57412 27257 57440
rect 27212 57400 27218 57412
rect 27341 57409 27353 57443
rect 27387 57440 27399 57443
rect 27798 57440 27804 57452
rect 27387 57412 27804 57440
rect 27387 57409 27399 57412
rect 27341 57403 27399 57409
rect 27798 57400 27804 57412
rect 27856 57400 27862 57452
rect 27893 57443 27951 57449
rect 27893 57409 27905 57443
rect 27939 57409 27951 57443
rect 27893 57403 27951 57409
rect 28905 57443 28963 57449
rect 28905 57409 28917 57443
rect 28951 57440 28963 57443
rect 29086 57440 29092 57452
rect 28951 57412 29092 57440
rect 28951 57409 28963 57412
rect 28905 57403 28963 57409
rect 24636 57344 26280 57372
rect 24636 57332 24642 57344
rect 26326 57332 26332 57384
rect 26384 57372 26390 57384
rect 27908 57372 27936 57403
rect 29086 57400 29092 57412
rect 29144 57400 29150 57452
rect 29472 57449 29500 57480
rect 29546 57468 29552 57520
rect 29604 57508 29610 57520
rect 41892 57517 41920 57548
rect 42150 57536 42156 57548
rect 42208 57576 42214 57588
rect 43346 57576 43352 57588
rect 42208 57548 43352 57576
rect 42208 57536 42214 57548
rect 43346 57536 43352 57548
rect 43404 57536 43410 57588
rect 36081 57511 36139 57517
rect 36081 57508 36093 57511
rect 29604 57480 31432 57508
rect 29604 57468 29610 57480
rect 29457 57443 29515 57449
rect 29457 57409 29469 57443
rect 29503 57440 29515 57443
rect 30374 57440 30380 57452
rect 29503 57412 30380 57440
rect 29503 57409 29515 57412
rect 29457 57403 29515 57409
rect 30374 57400 30380 57412
rect 30432 57400 30438 57452
rect 30834 57400 30840 57452
rect 30892 57440 30898 57452
rect 30929 57443 30987 57449
rect 30929 57440 30941 57443
rect 30892 57412 30941 57440
rect 30892 57400 30898 57412
rect 30929 57409 30941 57412
rect 30975 57409 30987 57443
rect 30929 57403 30987 57409
rect 26384 57344 27936 57372
rect 30285 57375 30343 57381
rect 26384 57332 26390 57344
rect 30285 57341 30297 57375
rect 30331 57372 30343 57375
rect 31294 57372 31300 57384
rect 30331 57344 31300 57372
rect 30331 57341 30343 57344
rect 30285 57335 30343 57341
rect 31294 57332 31300 57344
rect 31352 57332 31358 57384
rect 29178 57304 29184 57316
rect 23676 57276 23980 57304
rect 24044 57276 29184 57304
rect 20622 57196 20628 57248
rect 20680 57236 20686 57248
rect 23676 57236 23704 57276
rect 23842 57236 23848 57248
rect 20680 57208 23704 57236
rect 23803 57208 23848 57236
rect 20680 57196 20686 57208
rect 23842 57196 23848 57208
rect 23900 57196 23906 57248
rect 23952 57236 23980 57276
rect 29178 57264 29184 57276
rect 29236 57264 29242 57316
rect 29641 57307 29699 57313
rect 29641 57273 29653 57307
rect 29687 57304 29699 57307
rect 31404 57304 31432 57480
rect 32692 57480 36093 57508
rect 31754 57400 31760 57452
rect 31812 57440 31818 57452
rect 32692 57449 32720 57480
rect 36081 57477 36093 57480
rect 36127 57477 36139 57511
rect 36081 57471 36139 57477
rect 41877 57511 41935 57517
rect 41877 57477 41889 57511
rect 41923 57477 41935 57511
rect 41877 57471 41935 57477
rect 45554 57468 45560 57520
rect 45612 57508 45618 57520
rect 45833 57511 45891 57517
rect 45833 57508 45845 57511
rect 45612 57480 45845 57508
rect 45612 57468 45618 57480
rect 45833 57477 45845 57480
rect 45879 57477 45891 57511
rect 45833 57471 45891 57477
rect 45940 57480 50200 57508
rect 32677 57443 32735 57449
rect 32677 57440 32689 57443
rect 31812 57412 32689 57440
rect 31812 57400 31818 57412
rect 32677 57409 32689 57412
rect 32723 57409 32735 57443
rect 32677 57403 32735 57409
rect 32766 57400 32772 57452
rect 32824 57440 32830 57452
rect 33594 57440 33600 57452
rect 32824 57412 33600 57440
rect 32824 57400 32830 57412
rect 33594 57400 33600 57412
rect 33652 57440 33658 57452
rect 33965 57443 34023 57449
rect 33965 57440 33977 57443
rect 33652 57412 33977 57440
rect 33652 57400 33658 57412
rect 33965 57409 33977 57412
rect 34011 57409 34023 57443
rect 33965 57403 34023 57409
rect 34149 57443 34207 57449
rect 34149 57409 34161 57443
rect 34195 57409 34207 57443
rect 34149 57403 34207 57409
rect 32398 57372 32404 57384
rect 32359 57344 32404 57372
rect 32398 57332 32404 57344
rect 32456 57332 32462 57384
rect 32950 57332 32956 57384
rect 33008 57372 33014 57384
rect 34164 57372 34192 57403
rect 34238 57400 34244 57452
rect 34296 57440 34302 57452
rect 34296 57412 34341 57440
rect 34296 57400 34302 57412
rect 34514 57400 34520 57452
rect 34572 57440 34578 57452
rect 34698 57440 34704 57452
rect 34572 57412 34704 57440
rect 34572 57400 34578 57412
rect 34698 57400 34704 57412
rect 34756 57440 34762 57452
rect 34885 57443 34943 57449
rect 34885 57440 34897 57443
rect 34756 57412 34897 57440
rect 34756 57400 34762 57412
rect 34885 57409 34897 57412
rect 34931 57409 34943 57443
rect 35618 57440 35624 57452
rect 35579 57412 35624 57440
rect 34885 57403 34943 57409
rect 35618 57400 35624 57412
rect 35676 57440 35682 57452
rect 35802 57440 35808 57452
rect 35676 57412 35808 57440
rect 35676 57400 35682 57412
rect 35802 57400 35808 57412
rect 35860 57400 35866 57452
rect 35894 57400 35900 57452
rect 35952 57440 35958 57452
rect 36725 57443 36783 57449
rect 36725 57440 36737 57443
rect 35952 57412 36737 57440
rect 35952 57400 35958 57412
rect 36725 57409 36737 57412
rect 36771 57440 36783 57443
rect 37182 57440 37188 57452
rect 36771 57412 37188 57440
rect 36771 57409 36783 57412
rect 36725 57403 36783 57409
rect 37182 57400 37188 57412
rect 37240 57400 37246 57452
rect 37274 57400 37280 57452
rect 37332 57440 37338 57452
rect 38013 57443 38071 57449
rect 38013 57440 38025 57443
rect 37332 57412 38025 57440
rect 37332 57400 37338 57412
rect 38013 57409 38025 57412
rect 38059 57440 38071 57443
rect 38470 57440 38476 57452
rect 38059 57412 38476 57440
rect 38059 57409 38071 57412
rect 38013 57403 38071 57409
rect 38470 57400 38476 57412
rect 38528 57400 38534 57452
rect 40405 57443 40463 57449
rect 40405 57409 40417 57443
rect 40451 57440 40463 57443
rect 40678 57440 40684 57452
rect 40451 57412 40684 57440
rect 40451 57409 40463 57412
rect 40405 57403 40463 57409
rect 40678 57400 40684 57412
rect 40736 57400 40742 57452
rect 42061 57443 42119 57449
rect 42061 57409 42073 57443
rect 42107 57409 42119 57443
rect 42061 57403 42119 57409
rect 34330 57372 34336 57384
rect 33008 57344 33916 57372
rect 34164 57344 34336 57372
rect 33008 57332 33014 57344
rect 33781 57307 33839 57313
rect 33781 57304 33793 57307
rect 29687 57276 30696 57304
rect 31404 57276 33793 57304
rect 29687 57273 29699 57276
rect 29641 57267 29699 57273
rect 25682 57236 25688 57248
rect 23952 57208 25688 57236
rect 25682 57196 25688 57208
rect 25740 57196 25746 57248
rect 26697 57239 26755 57245
rect 26697 57205 26709 57239
rect 26743 57236 26755 57239
rect 27154 57236 27160 57248
rect 26743 57208 27160 57236
rect 26743 57205 26755 57208
rect 26697 57199 26755 57205
rect 27154 57196 27160 57208
rect 27212 57196 27218 57248
rect 27341 57239 27399 57245
rect 27341 57205 27353 57239
rect 27387 57236 27399 57239
rect 27430 57236 27436 57248
rect 27387 57208 27436 57236
rect 27387 57205 27399 57208
rect 27341 57199 27399 57205
rect 27430 57196 27436 57208
rect 27488 57196 27494 57248
rect 27522 57196 27528 57248
rect 27580 57236 27586 57248
rect 28810 57236 28816 57248
rect 27580 57208 28816 57236
rect 27580 57196 27586 57208
rect 28810 57196 28816 57208
rect 28868 57196 28874 57248
rect 30668 57236 30696 57276
rect 33781 57273 33793 57276
rect 33827 57273 33839 57307
rect 33888 57304 33916 57344
rect 34330 57332 34336 57344
rect 34388 57332 34394 57384
rect 34606 57332 34612 57384
rect 34664 57372 34670 57384
rect 37001 57375 37059 57381
rect 37001 57372 37013 57375
rect 34664 57344 37013 57372
rect 34664 57332 34670 57344
rect 37001 57341 37013 57344
rect 37047 57341 37059 57375
rect 37001 57335 37059 57341
rect 38289 57375 38347 57381
rect 38289 57341 38301 57375
rect 38335 57341 38347 57375
rect 40218 57372 40224 57384
rect 40179 57344 40224 57372
rect 38289 57335 38347 57341
rect 35437 57307 35495 57313
rect 35437 57304 35449 57307
rect 33888 57276 35449 57304
rect 33781 57267 33839 57273
rect 35437 57273 35449 57276
rect 35483 57273 35495 57307
rect 35437 57267 35495 57273
rect 33042 57236 33048 57248
rect 30668 57208 33048 57236
rect 33042 57196 33048 57208
rect 33100 57196 33106 57248
rect 33229 57239 33287 57245
rect 33229 57205 33241 57239
rect 33275 57236 33287 57239
rect 33318 57236 33324 57248
rect 33275 57208 33324 57236
rect 33275 57205 33287 57208
rect 33229 57199 33287 57205
rect 33318 57196 33324 57208
rect 33376 57236 33382 57248
rect 34238 57236 34244 57248
rect 33376 57208 34244 57236
rect 33376 57196 33382 57208
rect 34238 57196 34244 57208
rect 34296 57196 34302 57248
rect 34790 57236 34796 57248
rect 34751 57208 34796 57236
rect 34790 57196 34796 57208
rect 34848 57196 34854 57248
rect 35526 57196 35532 57248
rect 35584 57236 35590 57248
rect 38304 57236 38332 57335
rect 40218 57332 40224 57344
rect 40276 57332 40282 57384
rect 40313 57375 40371 57381
rect 40313 57341 40325 57375
rect 40359 57341 40371 57375
rect 40313 57335 40371 57341
rect 40328 57304 40356 57335
rect 40494 57332 40500 57384
rect 40552 57372 40558 57384
rect 42076 57372 42104 57403
rect 42794 57400 42800 57452
rect 42852 57440 42858 57452
rect 42889 57443 42947 57449
rect 42889 57440 42901 57443
rect 42852 57412 42901 57440
rect 42852 57400 42858 57412
rect 42889 57409 42901 57412
rect 42935 57440 42947 57443
rect 44082 57440 44088 57452
rect 42935 57412 44088 57440
rect 42935 57409 42947 57412
rect 42889 57403 42947 57409
rect 44082 57400 44088 57412
rect 44140 57400 44146 57452
rect 45462 57440 45468 57452
rect 44192 57412 45468 57440
rect 43070 57372 43076 57384
rect 40552 57344 40597 57372
rect 42076 57344 43076 57372
rect 40552 57332 40558 57344
rect 43070 57332 43076 57344
rect 43128 57372 43134 57384
rect 43165 57375 43223 57381
rect 43165 57372 43177 57375
rect 43128 57344 43177 57372
rect 43128 57332 43134 57344
rect 43165 57341 43177 57344
rect 43211 57341 43223 57375
rect 43165 57335 43223 57341
rect 43346 57332 43352 57384
rect 43404 57372 43410 57384
rect 44192 57372 44220 57412
rect 45462 57400 45468 57412
rect 45520 57440 45526 57452
rect 45940 57440 45968 57480
rect 45520 57412 45968 57440
rect 45520 57400 45526 57412
rect 46934 57400 46940 57452
rect 46992 57440 46998 57452
rect 47029 57443 47087 57449
rect 47029 57440 47041 57443
rect 46992 57412 47041 57440
rect 46992 57400 46998 57412
rect 47029 57409 47041 57412
rect 47075 57409 47087 57443
rect 47029 57403 47087 57409
rect 48314 57400 48320 57452
rect 48372 57440 48378 57452
rect 48501 57443 48559 57449
rect 48501 57440 48513 57443
rect 48372 57412 48513 57440
rect 48372 57400 48378 57412
rect 48501 57409 48513 57412
rect 48547 57409 48559 57443
rect 48501 57403 48559 57409
rect 49694 57400 49700 57452
rect 49752 57440 49758 57452
rect 49789 57443 49847 57449
rect 49789 57440 49801 57443
rect 49752 57412 49801 57440
rect 49752 57400 49758 57412
rect 49789 57409 49801 57412
rect 49835 57409 49847 57443
rect 49789 57403 49847 57409
rect 43404 57344 44220 57372
rect 43404 57332 43410 57344
rect 45002 57332 45008 57384
rect 45060 57372 45066 57384
rect 47305 57375 47363 57381
rect 47305 57372 47317 57375
rect 45060 57344 47317 57372
rect 45060 57332 45066 57344
rect 47305 57341 47317 57344
rect 47351 57341 47363 57375
rect 47305 57335 47363 57341
rect 47486 57332 47492 57384
rect 47544 57372 47550 57384
rect 48777 57375 48835 57381
rect 48777 57372 48789 57375
rect 47544 57344 48789 57372
rect 47544 57332 47550 57344
rect 48777 57341 48789 57344
rect 48823 57341 48835 57375
rect 48777 57335 48835 57341
rect 50065 57375 50123 57381
rect 50065 57341 50077 57375
rect 50111 57341 50123 57375
rect 50065 57335 50123 57341
rect 40236 57276 40356 57304
rect 40236 57248 40264 57276
rect 43990 57264 43996 57316
rect 44048 57304 44054 57316
rect 50080 57304 50108 57335
rect 44048 57276 50108 57304
rect 50172 57304 50200 57480
rect 52454 57468 52460 57520
rect 52512 57508 52518 57520
rect 52641 57511 52699 57517
rect 52641 57508 52653 57511
rect 52512 57480 52653 57508
rect 52512 57468 52518 57480
rect 52641 57477 52653 57480
rect 52687 57477 52699 57511
rect 52641 57471 52699 57477
rect 51074 57400 51080 57452
rect 51132 57440 51138 57452
rect 51445 57443 51503 57449
rect 51445 57440 51457 57443
rect 51132 57412 51457 57440
rect 51132 57400 51138 57412
rect 51445 57409 51457 57412
rect 51491 57409 51503 57443
rect 51445 57403 51503 57409
rect 52914 57400 52920 57452
rect 52972 57440 52978 57452
rect 53469 57443 53527 57449
rect 53469 57440 53481 57443
rect 52972 57412 53481 57440
rect 52972 57400 52978 57412
rect 53469 57409 53481 57412
rect 53515 57409 53527 57443
rect 53469 57403 53527 57409
rect 53834 57400 53840 57452
rect 53892 57440 53898 57452
rect 54202 57440 54208 57452
rect 53892 57412 54208 57440
rect 53892 57400 53898 57412
rect 54202 57400 54208 57412
rect 54260 57440 54266 57452
rect 54389 57443 54447 57449
rect 54389 57440 54401 57443
rect 54260 57412 54401 57440
rect 54260 57400 54266 57412
rect 54389 57409 54401 57412
rect 54435 57409 54447 57443
rect 54389 57403 54447 57409
rect 55214 57400 55220 57452
rect 55272 57440 55278 57452
rect 55585 57443 55643 57449
rect 55585 57440 55597 57443
rect 55272 57412 55597 57440
rect 55272 57400 55278 57412
rect 55585 57409 55597 57412
rect 55631 57409 55643 57443
rect 55585 57403 55643 57409
rect 55674 57400 55680 57452
rect 55732 57440 55738 57452
rect 56045 57443 56103 57449
rect 56045 57440 56057 57443
rect 55732 57412 56057 57440
rect 55732 57400 55738 57412
rect 56045 57409 56057 57412
rect 56091 57409 56103 57443
rect 56045 57403 56103 57409
rect 54573 57307 54631 57313
rect 54573 57304 54585 57307
rect 50172 57276 54585 57304
rect 44048 57264 44054 57276
rect 54573 57273 54585 57276
rect 54619 57273 54631 57307
rect 54573 57267 54631 57273
rect 35584 57208 38332 57236
rect 35584 57196 35590 57208
rect 40218 57196 40224 57248
rect 40276 57196 40282 57248
rect 41046 57236 41052 57248
rect 41007 57208 41052 57236
rect 41046 57196 41052 57208
rect 41104 57196 41110 57248
rect 41690 57236 41696 57248
rect 41651 57208 41696 57236
rect 41690 57196 41696 57208
rect 41748 57196 41754 57248
rect 44174 57236 44180 57248
rect 44135 57208 44180 57236
rect 44174 57196 44180 57208
rect 44232 57196 44238 57248
rect 44818 57236 44824 57248
rect 44779 57208 44824 57236
rect 44818 57196 44824 57208
rect 44876 57196 44882 57248
rect 44910 57196 44916 57248
rect 44968 57236 44974 57248
rect 45741 57239 45799 57245
rect 45741 57236 45753 57239
rect 44968 57208 45753 57236
rect 44968 57196 44974 57208
rect 45741 57205 45753 57208
rect 45787 57205 45799 57239
rect 46382 57236 46388 57248
rect 46343 57208 46388 57236
rect 45741 57199 45799 57205
rect 46382 57196 46388 57208
rect 46440 57196 46446 57248
rect 51626 57236 51632 57248
rect 51587 57208 51632 57236
rect 51626 57196 51632 57208
rect 51684 57196 51690 57248
rect 52730 57236 52736 57248
rect 52691 57208 52736 57236
rect 52730 57196 52736 57208
rect 52788 57196 52794 57248
rect 55398 57236 55404 57248
rect 55359 57208 55404 57236
rect 55398 57196 55404 57208
rect 55456 57196 55462 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 4614 56992 4620 57044
rect 4672 57032 4678 57044
rect 4709 57035 4767 57041
rect 4709 57032 4721 57035
rect 4672 57004 4721 57032
rect 4672 56992 4678 57004
rect 4709 57001 4721 57004
rect 4755 57001 4767 57035
rect 4709 56995 4767 57001
rect 10134 56992 10140 57044
rect 10192 57032 10198 57044
rect 10321 57035 10379 57041
rect 10321 57032 10333 57035
rect 10192 57004 10333 57032
rect 10192 56992 10198 57004
rect 10321 57001 10333 57004
rect 10367 57001 10379 57035
rect 10321 56995 10379 57001
rect 12894 56992 12900 57044
rect 12952 57032 12958 57044
rect 12989 57035 13047 57041
rect 12989 57032 13001 57035
rect 12952 57004 13001 57032
rect 12952 56992 12958 57004
rect 12989 57001 13001 57004
rect 13035 57001 13047 57035
rect 12989 56995 13047 57001
rect 15654 56992 15660 57044
rect 15712 57032 15718 57044
rect 16301 57035 16359 57041
rect 16301 57032 16313 57035
rect 15712 57004 16313 57032
rect 15712 56992 15718 57004
rect 16301 57001 16313 57004
rect 16347 57001 16359 57035
rect 16301 56995 16359 57001
rect 19889 57035 19947 57041
rect 19889 57001 19901 57035
rect 19935 57032 19947 57035
rect 19978 57032 19984 57044
rect 19935 57004 19984 57032
rect 19935 57001 19947 57004
rect 19889 56995 19947 57001
rect 19978 56992 19984 57004
rect 20036 56992 20042 57044
rect 21174 56992 21180 57044
rect 21232 57032 21238 57044
rect 21269 57035 21327 57041
rect 21269 57032 21281 57035
rect 21232 57004 21281 57032
rect 21232 56992 21238 57004
rect 21269 57001 21281 57004
rect 21315 57001 21327 57035
rect 23198 57032 23204 57044
rect 21269 56995 21327 57001
rect 22066 57004 23204 57032
rect 10962 56924 10968 56976
rect 11020 56964 11026 56976
rect 11149 56967 11207 56973
rect 11149 56964 11161 56967
rect 11020 56936 11161 56964
rect 11020 56924 11026 56936
rect 11149 56933 11161 56936
rect 11195 56964 11207 56967
rect 22066 56964 22094 57004
rect 23198 56992 23204 57004
rect 23256 56992 23262 57044
rect 23474 57032 23480 57044
rect 23387 57004 23480 57032
rect 23474 56992 23480 57004
rect 23532 57032 23538 57044
rect 24118 57032 24124 57044
rect 23532 57004 24124 57032
rect 23532 56992 23538 57004
rect 24118 56992 24124 57004
rect 24176 56992 24182 57044
rect 24578 57032 24584 57044
rect 24539 57004 24584 57032
rect 24578 56992 24584 57004
rect 24636 56992 24642 57044
rect 25038 57032 25044 57044
rect 24999 57004 25044 57032
rect 25038 56992 25044 57004
rect 25096 56992 25102 57044
rect 27798 56992 27804 57044
rect 27856 57032 27862 57044
rect 29086 57032 29092 57044
rect 27856 57004 28948 57032
rect 29047 57004 29092 57032
rect 27856 56992 27862 57004
rect 28920 56976 28948 57004
rect 29086 56992 29092 57004
rect 29144 56992 29150 57044
rect 29178 56992 29184 57044
rect 29236 57032 29242 57044
rect 30745 57035 30803 57041
rect 30745 57032 30757 57035
rect 29236 57004 30757 57032
rect 29236 56992 29242 57004
rect 30745 57001 30757 57004
rect 30791 57001 30803 57035
rect 30745 56995 30803 57001
rect 32674 56992 32680 57044
rect 32732 57032 32738 57044
rect 34241 57035 34299 57041
rect 34241 57032 34253 57035
rect 32732 57004 34253 57032
rect 32732 56992 32738 57004
rect 34241 57001 34253 57004
rect 34287 57001 34299 57035
rect 34241 56995 34299 57001
rect 40221 57035 40279 57041
rect 40221 57001 40233 57035
rect 40267 57032 40279 57035
rect 40494 57032 40500 57044
rect 40267 57004 40500 57032
rect 40267 57001 40279 57004
rect 40221 56995 40279 57001
rect 40494 56992 40500 57004
rect 40552 56992 40558 57044
rect 40770 56992 40776 57044
rect 40828 57032 40834 57044
rect 40828 57004 42656 57032
rect 40828 56992 40834 57004
rect 11195 56936 22094 56964
rect 22925 56967 22983 56973
rect 11195 56933 11207 56936
rect 11149 56927 11207 56933
rect 22925 56933 22937 56967
rect 22971 56964 22983 56967
rect 25314 56964 25320 56976
rect 22971 56936 25320 56964
rect 22971 56933 22983 56936
rect 22925 56927 22983 56933
rect 25314 56924 25320 56936
rect 25372 56924 25378 56976
rect 28166 56924 28172 56976
rect 28224 56964 28230 56976
rect 28353 56967 28411 56973
rect 28353 56964 28365 56967
rect 28224 56936 28365 56964
rect 28224 56924 28230 56936
rect 28353 56933 28365 56936
rect 28399 56933 28411 56967
rect 28902 56964 28908 56976
rect 28815 56936 28908 56964
rect 28353 56927 28411 56933
rect 28902 56924 28908 56936
rect 28960 56964 28966 56976
rect 32861 56967 32919 56973
rect 32861 56964 32873 56967
rect 28960 56936 29500 56964
rect 28960 56924 28966 56936
rect 16482 56856 16488 56908
rect 16540 56896 16546 56908
rect 26878 56896 26884 56908
rect 16540 56868 26884 56896
rect 16540 56856 16546 56868
rect 26878 56856 26884 56868
rect 26936 56856 26942 56908
rect 26970 56856 26976 56908
rect 27028 56896 27034 56908
rect 27617 56899 27675 56905
rect 27028 56868 27476 56896
rect 27028 56856 27034 56868
rect 23382 56828 23388 56840
rect 23343 56800 23388 56828
rect 23382 56788 23388 56800
rect 23440 56788 23446 56840
rect 23904 56831 23962 56837
rect 23904 56797 23916 56831
rect 23950 56828 23962 56831
rect 24026 56828 24032 56840
rect 23950 56800 24032 56828
rect 23950 56797 23962 56800
rect 23904 56791 23962 56797
rect 24026 56788 24032 56800
rect 24084 56788 24090 56840
rect 25222 56831 25280 56837
rect 25222 56797 25234 56831
rect 25268 56828 25280 56831
rect 25406 56828 25412 56840
rect 25268 56800 25412 56828
rect 25268 56797 25280 56800
rect 25222 56791 25280 56797
rect 25406 56788 25412 56800
rect 25464 56788 25470 56840
rect 25590 56828 25596 56840
rect 25551 56800 25596 56828
rect 25590 56788 25596 56800
rect 25648 56788 25654 56840
rect 25682 56788 25688 56840
rect 25740 56828 25746 56840
rect 26421 56831 26479 56837
rect 25740 56800 25785 56828
rect 25740 56788 25746 56800
rect 26421 56797 26433 56831
rect 26467 56828 26479 56831
rect 26510 56828 26516 56840
rect 26467 56800 26516 56828
rect 26467 56797 26479 56800
rect 26421 56791 26479 56797
rect 26510 56788 26516 56800
rect 26568 56788 26574 56840
rect 26602 56788 26608 56840
rect 26660 56828 26666 56840
rect 26660 56800 26705 56828
rect 26660 56788 26666 56800
rect 27062 56788 27068 56840
rect 27120 56828 27126 56840
rect 27448 56837 27476 56868
rect 27617 56865 27629 56899
rect 27663 56896 27675 56899
rect 29178 56896 29184 56908
rect 27663 56868 29184 56896
rect 27663 56865 27675 56868
rect 27617 56859 27675 56865
rect 29178 56856 29184 56868
rect 29236 56856 29242 56908
rect 27341 56831 27399 56837
rect 27341 56828 27353 56831
rect 27120 56800 27353 56828
rect 27120 56788 27126 56800
rect 27341 56797 27353 56800
rect 27387 56797 27399 56831
rect 27341 56791 27399 56797
rect 27433 56831 27491 56837
rect 27433 56797 27445 56831
rect 27479 56828 27491 56831
rect 27522 56828 27528 56840
rect 27479 56800 27528 56828
rect 27479 56797 27491 56800
rect 27433 56791 27491 56797
rect 27522 56788 27528 56800
rect 27580 56788 27586 56840
rect 27706 56828 27712 56840
rect 27667 56800 27712 56828
rect 27706 56788 27712 56800
rect 27764 56788 27770 56840
rect 28629 56831 28687 56837
rect 28276 56800 28580 56828
rect 27157 56763 27215 56769
rect 27157 56760 27169 56763
rect 6886 56732 27169 56760
rect 5442 56652 5448 56704
rect 5500 56692 5506 56704
rect 5629 56695 5687 56701
rect 5629 56692 5641 56695
rect 5500 56664 5641 56692
rect 5500 56652 5506 56664
rect 5629 56661 5641 56664
rect 5675 56692 5687 56695
rect 6886 56692 6914 56732
rect 27157 56729 27169 56732
rect 27203 56729 27215 56763
rect 27157 56723 27215 56729
rect 5675 56664 6914 56692
rect 5675 56661 5687 56664
rect 5629 56655 5687 56661
rect 23750 56652 23756 56704
rect 23808 56692 23814 56704
rect 23845 56695 23903 56701
rect 23845 56692 23857 56695
rect 23808 56664 23857 56692
rect 23808 56652 23814 56664
rect 23845 56661 23857 56664
rect 23891 56661 23903 56695
rect 23845 56655 23903 56661
rect 23934 56652 23940 56704
rect 23992 56692 23998 56704
rect 24029 56695 24087 56701
rect 24029 56692 24041 56695
rect 23992 56664 24041 56692
rect 23992 56652 23998 56664
rect 24029 56661 24041 56664
rect 24075 56661 24087 56695
rect 24029 56655 24087 56661
rect 25225 56695 25283 56701
rect 25225 56661 25237 56695
rect 25271 56692 25283 56695
rect 25498 56692 25504 56704
rect 25271 56664 25504 56692
rect 25271 56661 25283 56664
rect 25225 56655 25283 56661
rect 25498 56652 25504 56664
rect 25556 56652 25562 56704
rect 26237 56695 26295 56701
rect 26237 56661 26249 56695
rect 26283 56692 26295 56695
rect 26418 56692 26424 56704
rect 26283 56664 26424 56692
rect 26283 56661 26295 56664
rect 26237 56655 26295 56661
rect 26418 56652 26424 56664
rect 26476 56652 26482 56704
rect 27338 56652 27344 56704
rect 27396 56692 27402 56704
rect 28276 56692 28304 56800
rect 28350 56720 28356 56772
rect 28408 56760 28414 56772
rect 28552 56760 28580 56800
rect 28629 56797 28641 56831
rect 28675 56828 28687 56831
rect 28718 56828 28724 56840
rect 28675 56800 28724 56828
rect 28675 56797 28687 56800
rect 28629 56791 28687 56797
rect 28718 56788 28724 56800
rect 28776 56788 28782 56840
rect 28810 56788 28816 56840
rect 28868 56828 28874 56840
rect 29270 56828 29276 56840
rect 28868 56800 29276 56828
rect 28868 56788 28874 56800
rect 29270 56788 29276 56800
rect 29328 56788 29334 56840
rect 29472 56837 29500 56936
rect 29748 56936 32873 56964
rect 29546 56856 29552 56908
rect 29604 56896 29610 56908
rect 29604 56868 29649 56896
rect 29604 56856 29610 56868
rect 29457 56831 29515 56837
rect 29457 56797 29469 56831
rect 29503 56797 29515 56831
rect 29457 56791 29515 56797
rect 29641 56831 29699 56837
rect 29641 56797 29653 56831
rect 29687 56828 29699 56831
rect 29748 56828 29776 56936
rect 32861 56933 32873 56936
rect 32907 56933 32919 56967
rect 32861 56927 32919 56933
rect 33229 56967 33287 56973
rect 33229 56933 33241 56967
rect 33275 56964 33287 56967
rect 33318 56964 33324 56976
rect 33275 56936 33324 56964
rect 33275 56933 33287 56936
rect 33229 56927 33287 56933
rect 33318 56924 33324 56936
rect 33376 56924 33382 56976
rect 40310 56924 40316 56976
rect 40368 56964 40374 56976
rect 40589 56967 40647 56973
rect 40589 56964 40601 56967
rect 40368 56936 40601 56964
rect 40368 56924 40374 56936
rect 40589 56933 40601 56936
rect 40635 56933 40647 56967
rect 40589 56927 40647 56933
rect 41141 56967 41199 56973
rect 41141 56933 41153 56967
rect 41187 56933 41199 56967
rect 41141 56927 41199 56933
rect 30650 56856 30656 56908
rect 30708 56896 30714 56908
rect 31021 56899 31079 56905
rect 31021 56896 31033 56899
rect 30708 56868 31033 56896
rect 30708 56856 30714 56868
rect 31021 56865 31033 56868
rect 31067 56865 31079 56899
rect 31021 56859 31079 56865
rect 31110 56856 31116 56908
rect 31168 56896 31174 56908
rect 35345 56899 35403 56905
rect 31168 56868 32076 56896
rect 31168 56856 31174 56868
rect 29687 56800 29776 56828
rect 29687 56797 29699 56800
rect 29641 56791 29699 56797
rect 29656 56760 29684 56791
rect 29822 56788 29828 56840
rect 29880 56828 29886 56840
rect 30926 56828 30932 56840
rect 29880 56800 29925 56828
rect 30887 56800 30932 56828
rect 29880 56788 29886 56800
rect 30926 56788 30932 56800
rect 30984 56788 30990 56840
rect 31202 56788 31208 56840
rect 31260 56828 31266 56840
rect 31910 56831 31968 56837
rect 31260 56800 31305 56828
rect 31260 56788 31266 56800
rect 31910 56797 31922 56831
rect 31956 56828 31968 56831
rect 32048 56828 32076 56868
rect 35345 56865 35357 56899
rect 35391 56896 35403 56899
rect 35710 56896 35716 56908
rect 35391 56868 35716 56896
rect 35391 56865 35403 56868
rect 35345 56859 35403 56865
rect 35710 56856 35716 56868
rect 35768 56896 35774 56908
rect 37737 56899 37795 56905
rect 37737 56896 37749 56899
rect 35768 56868 37749 56896
rect 35768 56856 35774 56868
rect 37737 56865 37749 56868
rect 37783 56865 37795 56899
rect 37737 56859 37795 56865
rect 38013 56899 38071 56905
rect 38013 56865 38025 56899
rect 38059 56896 38071 56899
rect 38286 56896 38292 56908
rect 38059 56868 38292 56896
rect 38059 56865 38071 56868
rect 38013 56859 38071 56865
rect 38286 56856 38292 56868
rect 38344 56856 38350 56908
rect 40218 56896 40224 56908
rect 38626 56868 40224 56896
rect 32306 56828 32312 56840
rect 31956 56800 32076 56828
rect 32267 56800 32312 56828
rect 31956 56797 31968 56800
rect 31910 56791 31968 56797
rect 32306 56788 32312 56800
rect 32364 56788 32370 56840
rect 32401 56831 32459 56837
rect 32401 56797 32413 56831
rect 32447 56828 32459 56831
rect 32766 56828 32772 56840
rect 32447 56800 32772 56828
rect 32447 56797 32459 56800
rect 32401 56791 32459 56797
rect 32766 56788 32772 56800
rect 32824 56788 32830 56840
rect 33042 56788 33048 56840
rect 33100 56828 33106 56840
rect 33321 56831 33379 56837
rect 33100 56800 33145 56828
rect 33100 56788 33106 56800
rect 33321 56797 33333 56831
rect 33367 56828 33379 56831
rect 34330 56828 34336 56840
rect 33367 56800 34336 56828
rect 33367 56797 33379 56800
rect 33321 56791 33379 56797
rect 34330 56788 34336 56800
rect 34388 56788 34394 56840
rect 34514 56788 34520 56840
rect 34572 56828 34578 56840
rect 34885 56831 34943 56837
rect 34885 56828 34897 56831
rect 34572 56800 34897 56828
rect 34572 56788 34578 56800
rect 34885 56797 34897 56800
rect 34931 56828 34943 56831
rect 35066 56828 35072 56840
rect 34931 56800 35072 56828
rect 34931 56797 34943 56800
rect 34885 56791 34943 56797
rect 35066 56788 35072 56800
rect 35124 56788 35130 56840
rect 35253 56831 35311 56837
rect 35253 56797 35265 56831
rect 35299 56828 35311 56831
rect 35526 56828 35532 56840
rect 35299 56800 35532 56828
rect 35299 56797 35311 56800
rect 35253 56791 35311 56797
rect 35526 56788 35532 56800
rect 35584 56788 35590 56840
rect 35989 56831 36047 56837
rect 35989 56828 36001 56831
rect 35636 56800 36001 56828
rect 35158 56760 35164 56772
rect 28408 56732 28453 56760
rect 28552 56732 29684 56760
rect 29748 56732 32352 56760
rect 28408 56720 28414 56732
rect 28534 56692 28540 56704
rect 27396 56664 28304 56692
rect 28495 56664 28540 56692
rect 27396 56652 27402 56664
rect 28534 56652 28540 56664
rect 28592 56652 28598 56704
rect 29178 56652 29184 56704
rect 29236 56692 29242 56704
rect 29748 56692 29776 56732
rect 29236 56664 29776 56692
rect 29236 56652 29242 56664
rect 31754 56652 31760 56704
rect 31812 56692 31818 56704
rect 31812 56664 31857 56692
rect 31812 56652 31818 56664
rect 31938 56652 31944 56704
rect 31996 56692 32002 56704
rect 32324 56692 32352 56732
rect 33060 56732 35164 56760
rect 33060 56692 33088 56732
rect 35158 56720 35164 56732
rect 35216 56720 35222 56772
rect 31996 56664 32041 56692
rect 32324 56664 33088 56692
rect 31996 56652 32002 56664
rect 33686 56652 33692 56704
rect 33744 56692 33750 56704
rect 34977 56695 35035 56701
rect 34977 56692 34989 56695
rect 33744 56664 34989 56692
rect 33744 56652 33750 56664
rect 34977 56661 34989 56664
rect 35023 56661 35035 56695
rect 34977 56655 35035 56661
rect 35066 56652 35072 56704
rect 35124 56692 35130 56704
rect 35636 56692 35664 56800
rect 35989 56797 36001 56800
rect 36035 56797 36047 56831
rect 35989 56791 36047 56797
rect 36265 56831 36323 56837
rect 36265 56797 36277 56831
rect 36311 56797 36323 56831
rect 36446 56828 36452 56840
rect 36407 56800 36452 56828
rect 36265 56791 36323 56797
rect 36280 56760 36308 56791
rect 36446 56788 36452 56800
rect 36504 56788 36510 56840
rect 36722 56828 36728 56840
rect 36683 56800 36728 56828
rect 36722 56788 36728 56800
rect 36780 56788 36786 56840
rect 37918 56828 37924 56840
rect 37879 56800 37924 56828
rect 37918 56788 37924 56800
rect 37976 56788 37982 56840
rect 38102 56828 38108 56840
rect 38063 56800 38108 56828
rect 38102 56788 38108 56800
rect 38160 56788 38166 56840
rect 38197 56831 38255 56837
rect 38197 56797 38209 56831
rect 38243 56828 38255 56831
rect 38626 56828 38654 56868
rect 40218 56856 40224 56868
rect 40276 56856 40282 56908
rect 41156 56896 41184 56927
rect 40420 56868 41184 56896
rect 38243 56800 38654 56828
rect 38243 56797 38255 56800
rect 38197 56791 38255 56797
rect 38746 56788 38752 56840
rect 38804 56828 38810 56840
rect 40420 56837 40448 56868
rect 41598 56856 41604 56908
rect 41656 56896 41662 56908
rect 41785 56899 41843 56905
rect 41785 56896 41797 56899
rect 41656 56868 41797 56896
rect 41656 56856 41662 56868
rect 41785 56865 41797 56868
rect 41831 56865 41843 56899
rect 41785 56859 41843 56865
rect 40405 56831 40463 56837
rect 38804 56800 38849 56828
rect 38804 56788 38810 56800
rect 40405 56797 40417 56831
rect 40451 56797 40463 56831
rect 40678 56828 40684 56840
rect 40639 56800 40684 56828
rect 40405 56791 40463 56797
rect 40678 56788 40684 56800
rect 40736 56788 40742 56840
rect 41322 56804 41328 56856
rect 41380 56804 41386 56856
rect 41693 56831 41751 56837
rect 41322 56797 41334 56804
rect 41368 56797 41380 56804
rect 41322 56791 41380 56797
rect 41693 56797 41705 56831
rect 41739 56828 41751 56831
rect 42150 56828 42156 56840
rect 41739 56800 42156 56828
rect 41739 56797 41751 56800
rect 41693 56791 41751 56797
rect 42150 56788 42156 56800
rect 42208 56788 42214 56840
rect 42628 56828 42656 57004
rect 47394 56992 47400 57044
rect 47452 57032 47458 57044
rect 48133 57035 48191 57041
rect 48133 57032 48145 57035
rect 47452 57004 48145 57032
rect 47452 56992 47458 57004
rect 48133 57001 48145 57004
rect 48179 57001 48191 57035
rect 48133 56995 48191 57001
rect 48774 56992 48780 57044
rect 48832 57032 48838 57044
rect 49421 57035 49479 57041
rect 49421 57032 49433 57035
rect 48832 57004 49433 57032
rect 48832 56992 48838 57004
rect 49421 57001 49433 57004
rect 49467 57001 49479 57035
rect 49421 56995 49479 57001
rect 50154 56992 50160 57044
rect 50212 57032 50218 57044
rect 50709 57035 50767 57041
rect 50709 57032 50721 57035
rect 50212 57004 50721 57032
rect 50212 56992 50218 57004
rect 50709 57001 50721 57004
rect 50755 57001 50767 57035
rect 50709 56995 50767 57001
rect 51534 56992 51540 57044
rect 51592 57032 51598 57044
rect 52181 57035 52239 57041
rect 52181 57032 52193 57035
rect 51592 57004 52193 57032
rect 51592 56992 51598 57004
rect 52181 57001 52193 57004
rect 52227 57001 52239 57035
rect 52181 56995 52239 57001
rect 53374 56992 53380 57044
rect 53432 57032 53438 57044
rect 53469 57035 53527 57041
rect 53469 57032 53481 57035
rect 53432 57004 53481 57032
rect 53432 56992 53438 57004
rect 53469 57001 53481 57004
rect 53515 57001 53527 57035
rect 53469 56995 53527 57001
rect 54294 56992 54300 57044
rect 54352 57032 54358 57044
rect 54389 57035 54447 57041
rect 54389 57032 54401 57035
rect 54352 57004 54401 57032
rect 54352 56992 54358 57004
rect 54389 57001 54401 57004
rect 54435 57001 54447 57035
rect 54389 56995 54447 57001
rect 54754 56992 54760 57044
rect 54812 57032 54818 57044
rect 55033 57035 55091 57041
rect 55033 57032 55045 57035
rect 54812 57004 55045 57032
rect 54812 56992 54818 57004
rect 55033 57001 55045 57004
rect 55079 57001 55091 57035
rect 55033 56995 55091 57001
rect 55214 56992 55220 57044
rect 55272 57032 55278 57044
rect 55677 57035 55735 57041
rect 55677 57032 55689 57035
rect 55272 57004 55689 57032
rect 55272 56992 55278 57004
rect 55677 57001 55689 57004
rect 55723 57001 55735 57035
rect 55677 56995 55735 57001
rect 56134 56992 56140 57044
rect 56192 57032 56198 57044
rect 56229 57035 56287 57041
rect 56229 57032 56241 57035
rect 56192 57004 56241 57032
rect 56192 56992 56198 57004
rect 56229 57001 56241 57004
rect 56275 57001 56287 57035
rect 56229 56995 56287 57001
rect 43806 56964 43812 56976
rect 43767 56936 43812 56964
rect 43806 56924 43812 56936
rect 43864 56924 43870 56976
rect 45462 56964 45468 56976
rect 44652 56936 45468 56964
rect 42797 56899 42855 56905
rect 42797 56865 42809 56899
rect 42843 56896 42855 56899
rect 43717 56899 43775 56905
rect 43717 56896 43729 56899
rect 42843 56868 43729 56896
rect 42843 56865 42855 56868
rect 42797 56859 42855 56865
rect 43717 56865 43729 56868
rect 43763 56865 43775 56899
rect 43898 56896 43904 56908
rect 43859 56868 43904 56896
rect 43717 56859 43775 56865
rect 43898 56856 43904 56868
rect 43956 56856 43962 56908
rect 42981 56831 43039 56837
rect 42981 56828 42993 56831
rect 42628 56800 42993 56828
rect 42981 56797 42993 56800
rect 43027 56797 43039 56831
rect 43162 56828 43168 56840
rect 43123 56800 43168 56828
rect 42981 56791 43039 56797
rect 36538 56760 36544 56772
rect 36280 56732 36544 56760
rect 36538 56720 36544 56732
rect 36596 56760 36602 56772
rect 41506 56760 41512 56772
rect 36596 56732 41512 56760
rect 36596 56720 36602 56732
rect 41506 56720 41512 56732
rect 41564 56720 41570 56772
rect 42996 56760 43024 56791
rect 43162 56788 43168 56800
rect 43220 56788 43226 56840
rect 43257 56831 43315 56837
rect 43257 56797 43269 56831
rect 43303 56828 43315 56831
rect 43990 56828 43996 56840
rect 43303 56800 43996 56828
rect 43303 56797 43315 56800
rect 43257 56791 43315 56797
rect 43990 56788 43996 56800
rect 44048 56828 44054 56840
rect 44177 56831 44235 56837
rect 44177 56828 44189 56831
rect 44048 56800 44189 56828
rect 44048 56788 44054 56800
rect 44177 56797 44189 56800
rect 44223 56797 44235 56831
rect 44177 56791 44235 56797
rect 44545 56831 44603 56837
rect 44545 56797 44557 56831
rect 44591 56828 44603 56831
rect 44652 56828 44680 56936
rect 45462 56924 45468 56936
rect 45520 56924 45526 56976
rect 46014 56924 46020 56976
rect 46072 56964 46078 56976
rect 47489 56967 47547 56973
rect 47489 56964 47501 56967
rect 46072 56936 47501 56964
rect 46072 56924 46078 56936
rect 47489 56933 47501 56936
rect 47535 56933 47547 56967
rect 47489 56927 47547 56933
rect 49234 56924 49240 56976
rect 49292 56964 49298 56976
rect 50065 56967 50123 56973
rect 50065 56964 50077 56967
rect 49292 56936 50077 56964
rect 49292 56924 49298 56936
rect 50065 56933 50077 56936
rect 50111 56933 50123 56967
rect 50065 56927 50123 56933
rect 50614 56924 50620 56976
rect 50672 56964 50678 56976
rect 51353 56967 51411 56973
rect 51353 56964 51365 56967
rect 50672 56936 51365 56964
rect 50672 56924 50678 56936
rect 51353 56933 51365 56936
rect 51399 56933 51411 56967
rect 51353 56927 51411 56933
rect 51994 56924 52000 56976
rect 52052 56964 52058 56976
rect 52825 56967 52883 56973
rect 52825 56964 52837 56967
rect 52052 56936 52837 56964
rect 52052 56924 52058 56936
rect 52825 56933 52837 56936
rect 52871 56933 52883 56967
rect 52825 56927 52883 56933
rect 47854 56856 47860 56908
rect 47912 56896 47918 56908
rect 48777 56899 48835 56905
rect 48777 56896 48789 56899
rect 47912 56868 48789 56896
rect 47912 56856 47918 56868
rect 48777 56865 48789 56868
rect 48823 56865 48835 56899
rect 48777 56859 48835 56865
rect 45186 56828 45192 56840
rect 44591 56800 44680 56828
rect 45147 56800 45192 56828
rect 44591 56797 44603 56800
rect 44545 56791 44603 56797
rect 45186 56788 45192 56800
rect 45244 56788 45250 56840
rect 46198 56828 46204 56840
rect 46159 56800 46204 56828
rect 46198 56788 46204 56800
rect 46256 56788 46262 56840
rect 46750 56788 46756 56840
rect 46808 56828 46814 56840
rect 47029 56831 47087 56837
rect 47029 56828 47041 56831
rect 46808 56800 47041 56828
rect 46808 56788 46814 56800
rect 47029 56797 47041 56800
rect 47075 56797 47087 56831
rect 47029 56791 47087 56797
rect 42996 56732 46888 56760
rect 36078 56692 36084 56704
rect 35124 56664 35664 56692
rect 36039 56664 36084 56692
rect 35124 56652 35130 56664
rect 36078 56652 36084 56664
rect 36136 56652 36142 56704
rect 36170 56652 36176 56704
rect 36228 56692 36234 56704
rect 38979 56695 39037 56701
rect 38979 56692 38991 56695
rect 36228 56664 38991 56692
rect 36228 56652 36234 56664
rect 38979 56661 38991 56664
rect 39025 56661 39037 56695
rect 38979 56655 39037 56661
rect 40310 56652 40316 56704
rect 40368 56692 40374 56704
rect 41325 56695 41383 56701
rect 41325 56692 41337 56695
rect 40368 56664 41337 56692
rect 40368 56652 40374 56664
rect 41325 56661 41337 56664
rect 41371 56661 41383 56695
rect 41325 56655 41383 56661
rect 41414 56652 41420 56704
rect 41472 56692 41478 56704
rect 42337 56695 42395 56701
rect 42337 56692 42349 56695
rect 41472 56664 42349 56692
rect 41472 56652 41478 56664
rect 42337 56661 42349 56664
rect 42383 56692 42395 56695
rect 42426 56692 42432 56704
rect 42383 56664 42432 56692
rect 42383 56661 42395 56664
rect 42337 56655 42395 56661
rect 42426 56652 42432 56664
rect 42484 56652 42490 56704
rect 42610 56652 42616 56704
rect 42668 56692 42674 56704
rect 46860 56701 46888 56732
rect 45005 56695 45063 56701
rect 45005 56692 45017 56695
rect 42668 56664 45017 56692
rect 42668 56652 42674 56664
rect 45005 56661 45017 56664
rect 45051 56661 45063 56695
rect 45005 56655 45063 56661
rect 46845 56695 46903 56701
rect 46845 56661 46857 56695
rect 46891 56661 46903 56695
rect 46845 56655 46903 56661
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 23474 56488 23480 56500
rect 23435 56460 23480 56488
rect 23474 56448 23480 56460
rect 23532 56448 23538 56500
rect 26510 56448 26516 56500
rect 26568 56488 26574 56500
rect 26697 56491 26755 56497
rect 26697 56488 26709 56491
rect 26568 56460 26709 56488
rect 26568 56448 26574 56460
rect 26697 56457 26709 56460
rect 26743 56457 26755 56491
rect 26878 56488 26884 56500
rect 26839 56460 26884 56488
rect 26697 56451 26755 56457
rect 17862 56380 17868 56432
rect 17920 56420 17926 56432
rect 26712 56420 26740 56451
rect 26878 56448 26884 56460
rect 26936 56448 26942 56500
rect 27706 56448 27712 56500
rect 27764 56488 27770 56500
rect 27985 56491 28043 56497
rect 27985 56488 27997 56491
rect 27764 56460 27997 56488
rect 27764 56448 27770 56460
rect 27985 56457 27997 56460
rect 28031 56457 28043 56491
rect 27985 56451 28043 56457
rect 28258 56448 28264 56500
rect 28316 56488 28322 56500
rect 29822 56488 29828 56500
rect 28316 56460 29828 56488
rect 28316 56448 28322 56460
rect 29822 56448 29828 56460
rect 29880 56448 29886 56500
rect 31202 56448 31208 56500
rect 31260 56488 31266 56500
rect 31481 56491 31539 56497
rect 31481 56488 31493 56491
rect 31260 56460 31493 56488
rect 31260 56448 31266 56460
rect 31481 56457 31493 56460
rect 31527 56457 31539 56491
rect 34790 56488 34796 56500
rect 31481 56451 31539 56457
rect 33152 56460 34796 56488
rect 26970 56420 26976 56432
rect 17920 56392 26372 56420
rect 26712 56392 26976 56420
rect 17920 56380 17926 56392
rect 22554 56312 22560 56364
rect 22612 56352 22618 56364
rect 22649 56355 22707 56361
rect 22649 56352 22661 56355
rect 22612 56324 22661 56352
rect 22612 56312 22618 56324
rect 22649 56321 22661 56324
rect 22695 56321 22707 56355
rect 22649 56315 22707 56321
rect 23293 56355 23351 56361
rect 23293 56321 23305 56355
rect 23339 56352 23351 56355
rect 23842 56352 23848 56364
rect 23339 56324 23848 56352
rect 23339 56321 23351 56324
rect 23293 56315 23351 56321
rect 23842 56312 23848 56324
rect 23900 56312 23906 56364
rect 23937 56355 23995 56361
rect 23937 56321 23949 56355
rect 23983 56321 23995 56355
rect 25498 56352 25504 56364
rect 25459 56324 25504 56352
rect 23937 56315 23995 56321
rect 23952 56284 23980 56315
rect 25498 56312 25504 56324
rect 25556 56312 25562 56364
rect 26234 56352 26240 56364
rect 26195 56324 26240 56352
rect 26234 56312 26240 56324
rect 26292 56312 26298 56364
rect 22112 56256 23980 56284
rect 5350 56108 5356 56160
rect 5408 56148 5414 56160
rect 22112 56157 22140 56256
rect 23952 56216 23980 56256
rect 24213 56287 24271 56293
rect 24213 56253 24225 56287
rect 24259 56284 24271 56287
rect 24302 56284 24308 56296
rect 24259 56256 24308 56284
rect 24259 56253 24271 56256
rect 24213 56247 24271 56253
rect 24302 56244 24308 56256
rect 24360 56284 24366 56296
rect 24762 56284 24768 56296
rect 24360 56256 24768 56284
rect 24360 56244 24366 56256
rect 24762 56244 24768 56256
rect 24820 56284 24826 56296
rect 25317 56287 25375 56293
rect 25317 56284 25329 56287
rect 24820 56256 25329 56284
rect 24820 56244 24826 56256
rect 25317 56253 25329 56256
rect 25363 56253 25375 56287
rect 26344 56284 26372 56392
rect 26970 56380 26976 56392
rect 27028 56380 27034 56432
rect 27430 56380 27436 56432
rect 27488 56420 27494 56432
rect 27488 56392 29132 56420
rect 27488 56380 27494 56392
rect 26756 56355 26814 56361
rect 26756 56321 26768 56355
rect 26802 56352 26814 56355
rect 26878 56352 26884 56364
rect 26802 56324 26884 56352
rect 26802 56321 26814 56324
rect 26756 56315 26814 56321
rect 26878 56312 26884 56324
rect 26936 56312 26942 56364
rect 27338 56352 27344 56364
rect 27299 56324 27344 56352
rect 27338 56312 27344 56324
rect 27396 56312 27402 56364
rect 27525 56355 27583 56361
rect 27525 56321 27537 56355
rect 27571 56352 27583 56355
rect 27614 56352 27620 56364
rect 27571 56324 27620 56352
rect 27571 56321 27583 56324
rect 27525 56315 27583 56321
rect 27614 56312 27620 56324
rect 27672 56312 27678 56364
rect 27706 56312 27712 56364
rect 27764 56352 27770 56364
rect 28166 56352 28172 56364
rect 27764 56324 28172 56352
rect 27764 56312 27770 56324
rect 28166 56312 28172 56324
rect 28224 56312 28230 56364
rect 28353 56355 28411 56361
rect 28353 56321 28365 56355
rect 28399 56352 28411 56355
rect 28442 56352 28448 56364
rect 28399 56324 28448 56352
rect 28399 56321 28411 56324
rect 28353 56315 28411 56321
rect 28442 56312 28448 56324
rect 28500 56312 28506 56364
rect 29104 56361 29132 56392
rect 29270 56380 29276 56432
rect 29328 56420 29334 56432
rect 29328 56392 29592 56420
rect 29328 56380 29334 56392
rect 29089 56355 29147 56361
rect 29089 56321 29101 56355
rect 29135 56321 29147 56355
rect 29089 56315 29147 56321
rect 29178 56312 29184 56364
rect 29236 56352 29242 56364
rect 29564 56361 29592 56392
rect 30098 56380 30104 56432
rect 30156 56420 30162 56432
rect 32950 56420 32956 56432
rect 30156 56392 32956 56420
rect 30156 56380 30162 56392
rect 32950 56380 32956 56392
rect 33008 56380 33014 56432
rect 29365 56355 29423 56361
rect 29365 56352 29377 56355
rect 29236 56324 29377 56352
rect 29236 56312 29242 56324
rect 29365 56321 29377 56324
rect 29411 56321 29423 56355
rect 29365 56315 29423 56321
rect 29549 56355 29607 56361
rect 29549 56321 29561 56355
rect 29595 56321 29607 56355
rect 29549 56315 29607 56321
rect 29914 56312 29920 56364
rect 29972 56352 29978 56364
rect 30009 56355 30067 56361
rect 30009 56352 30021 56355
rect 29972 56324 30021 56352
rect 29972 56312 29978 56324
rect 30009 56321 30021 56324
rect 30055 56321 30067 56355
rect 30009 56315 30067 56321
rect 31665 56355 31723 56361
rect 31665 56321 31677 56355
rect 31711 56352 31723 56355
rect 31754 56352 31760 56364
rect 31711 56324 31760 56352
rect 31711 56321 31723 56324
rect 31665 56315 31723 56321
rect 31754 56312 31760 56324
rect 31812 56312 31818 56364
rect 32214 56312 32220 56364
rect 32272 56352 32278 56364
rect 32401 56355 32459 56361
rect 32401 56352 32413 56355
rect 32272 56324 32413 56352
rect 32272 56312 32278 56324
rect 32401 56321 32413 56324
rect 32447 56321 32459 56355
rect 33152 56352 33180 56460
rect 34790 56448 34796 56460
rect 34848 56448 34854 56500
rect 35158 56448 35164 56500
rect 35216 56488 35222 56500
rect 35345 56491 35403 56497
rect 35345 56488 35357 56491
rect 35216 56460 35357 56488
rect 35216 56448 35222 56460
rect 35345 56457 35357 56460
rect 35391 56457 35403 56491
rect 35345 56451 35403 56457
rect 36446 56448 36452 56500
rect 36504 56488 36510 56500
rect 36504 56460 36676 56488
rect 36504 56448 36510 56460
rect 35710 56420 35716 56432
rect 33428 56392 34652 56420
rect 35671 56392 35716 56420
rect 33318 56352 33324 56364
rect 32401 56315 32459 56321
rect 33060 56324 33180 56352
rect 33279 56324 33324 56352
rect 28905 56287 28963 56293
rect 28905 56284 28917 56287
rect 26344 56256 28917 56284
rect 25317 56247 25375 56253
rect 28905 56253 28917 56256
rect 28951 56253 28963 56287
rect 28905 56247 28963 56253
rect 29273 56287 29331 56293
rect 29273 56253 29285 56287
rect 29319 56253 29331 56287
rect 29273 56247 29331 56253
rect 26326 56216 26332 56228
rect 23952 56188 26188 56216
rect 26287 56188 26332 56216
rect 22097 56151 22155 56157
rect 22097 56148 22109 56151
rect 5408 56120 22109 56148
rect 5408 56108 5414 56120
rect 22097 56117 22109 56120
rect 22143 56117 22155 56151
rect 25682 56148 25688 56160
rect 25643 56120 25688 56148
rect 22097 56111 22155 56117
rect 25682 56108 25688 56120
rect 25740 56108 25746 56160
rect 26160 56148 26188 56188
rect 26326 56176 26332 56188
rect 26384 56176 26390 56228
rect 27525 56219 27583 56225
rect 27525 56185 27537 56219
rect 27571 56216 27583 56219
rect 29181 56219 29239 56225
rect 29181 56216 29193 56219
rect 27571 56188 29193 56216
rect 27571 56185 27583 56188
rect 27525 56179 27583 56185
rect 29181 56185 29193 56188
rect 29227 56185 29239 56219
rect 29288 56216 29316 56247
rect 31110 56244 31116 56296
rect 31168 56284 31174 56296
rect 31570 56284 31576 56296
rect 31168 56256 31576 56284
rect 31168 56244 31174 56256
rect 31570 56244 31576 56256
rect 31628 56284 31634 56296
rect 31941 56287 31999 56293
rect 31941 56284 31953 56287
rect 31628 56256 31953 56284
rect 31628 56244 31634 56256
rect 31941 56253 31953 56256
rect 31987 56284 31999 56287
rect 33060 56284 33088 56324
rect 33318 56312 33324 56324
rect 33376 56312 33382 56364
rect 33428 56361 33456 56392
rect 34624 56364 34652 56392
rect 35710 56380 35716 56392
rect 35768 56380 35774 56432
rect 36648 56429 36676 56460
rect 36814 56448 36820 56500
rect 36872 56488 36878 56500
rect 41046 56488 41052 56500
rect 36872 56460 41052 56488
rect 36872 56448 36878 56460
rect 41046 56448 41052 56460
rect 41104 56448 41110 56500
rect 43254 56448 43260 56500
rect 43312 56488 43318 56500
rect 46382 56488 46388 56500
rect 43312 56460 46388 56488
rect 43312 56448 43318 56460
rect 46382 56448 46388 56460
rect 46440 56448 46446 56500
rect 48314 56488 48320 56500
rect 48275 56460 48320 56488
rect 48314 56448 48320 56460
rect 48372 56448 48378 56500
rect 49694 56488 49700 56500
rect 49655 56460 49700 56488
rect 49694 56448 49700 56460
rect 49752 56448 49758 56500
rect 51074 56448 51080 56500
rect 51132 56488 51138 56500
rect 51261 56491 51319 56497
rect 51261 56488 51273 56491
rect 51132 56460 51273 56488
rect 51132 56448 51138 56460
rect 51261 56457 51273 56460
rect 51307 56457 51319 56491
rect 52454 56488 52460 56500
rect 52415 56460 52460 56488
rect 51261 56451 51319 56457
rect 52454 56448 52460 56460
rect 52512 56448 52518 56500
rect 54202 56488 54208 56500
rect 54163 56460 54208 56488
rect 54202 56448 54208 56460
rect 54260 56448 54266 56500
rect 36633 56423 36691 56429
rect 36633 56389 36645 56423
rect 36679 56420 36691 56423
rect 39022 56420 39028 56432
rect 36679 56392 39028 56420
rect 36679 56389 36691 56392
rect 36633 56383 36691 56389
rect 39022 56380 39028 56392
rect 39080 56380 39086 56432
rect 41690 56420 41696 56432
rect 40052 56392 41696 56420
rect 33413 56355 33471 56361
rect 33413 56321 33425 56355
rect 33459 56321 33471 56355
rect 33594 56352 33600 56364
rect 33555 56324 33600 56352
rect 33413 56315 33471 56321
rect 33594 56312 33600 56324
rect 33652 56312 33658 56364
rect 33689 56355 33747 56361
rect 33689 56321 33701 56355
rect 33735 56352 33747 56355
rect 34149 56355 34207 56361
rect 34149 56352 34161 56355
rect 33735 56324 34161 56352
rect 33735 56321 33747 56324
rect 33689 56315 33747 56321
rect 34149 56321 34161 56324
rect 34195 56321 34207 56355
rect 34149 56315 34207 56321
rect 34333 56355 34391 56361
rect 34333 56321 34345 56355
rect 34379 56321 34391 56355
rect 34606 56352 34612 56364
rect 34567 56324 34612 56352
rect 34333 56315 34391 56321
rect 31987 56256 33088 56284
rect 31987 56253 31999 56256
rect 31941 56247 31999 56253
rect 33134 56244 33140 56296
rect 33192 56284 33198 56296
rect 34348 56284 34376 56315
rect 34606 56312 34612 56324
rect 34664 56312 34670 56364
rect 35526 56352 35532 56364
rect 35487 56324 35532 56352
rect 35526 56312 35532 56324
rect 35584 56312 35590 56364
rect 36449 56355 36507 56361
rect 36449 56321 36461 56355
rect 36495 56352 36507 56355
rect 36538 56352 36544 56364
rect 36495 56324 36544 56352
rect 36495 56321 36507 56324
rect 36449 56315 36507 56321
rect 36538 56312 36544 56324
rect 36596 56312 36602 56364
rect 36722 56312 36728 56364
rect 36780 56352 36786 56364
rect 40052 56361 40080 56392
rect 41690 56380 41696 56392
rect 41748 56380 41754 56432
rect 43162 56380 43168 56432
rect 43220 56420 43226 56432
rect 43346 56420 43352 56432
rect 43220 56392 43352 56420
rect 43220 56380 43226 56392
rect 43346 56380 43352 56392
rect 43404 56380 43410 56432
rect 43714 56380 43720 56432
rect 43772 56420 43778 56432
rect 46198 56420 46204 56432
rect 43772 56392 46204 56420
rect 43772 56380 43778 56392
rect 46198 56380 46204 56392
rect 46256 56380 46262 56432
rect 38749 56355 38807 56361
rect 36780 56324 36825 56352
rect 36780 56312 36786 56324
rect 38749 56321 38761 56355
rect 38795 56321 38807 56355
rect 38749 56315 38807 56321
rect 40037 56355 40095 56361
rect 40037 56321 40049 56355
rect 40083 56321 40095 56355
rect 40037 56315 40095 56321
rect 40129 56355 40187 56361
rect 40129 56321 40141 56355
rect 40175 56321 40187 56355
rect 40129 56315 40187 56321
rect 33192 56256 34376 56284
rect 38105 56287 38163 56293
rect 33192 56244 33198 56256
rect 38105 56253 38117 56287
rect 38151 56284 38163 56287
rect 38562 56284 38568 56296
rect 38151 56256 38568 56284
rect 38151 56253 38163 56256
rect 38105 56247 38163 56253
rect 38562 56244 38568 56256
rect 38620 56244 38626 56296
rect 36265 56219 36323 56225
rect 36265 56216 36277 56219
rect 29288 56188 36277 56216
rect 29181 56179 29239 56185
rect 36265 56185 36277 56188
rect 36311 56185 36323 56219
rect 36265 56179 36323 56185
rect 37829 56219 37887 56225
rect 37829 56185 37841 56219
rect 37875 56216 37887 56219
rect 38286 56216 38292 56228
rect 37875 56188 38292 56216
rect 37875 56185 37887 56188
rect 37829 56179 37887 56185
rect 38286 56176 38292 56188
rect 38344 56176 38350 56228
rect 38764 56216 38792 56315
rect 38930 56284 38936 56296
rect 38891 56256 38936 56284
rect 38930 56244 38936 56256
rect 38988 56244 38994 56296
rect 40144 56216 40172 56315
rect 40218 56312 40224 56364
rect 40276 56352 40282 56364
rect 40359 56355 40417 56361
rect 40276 56324 40321 56352
rect 40276 56312 40282 56324
rect 40359 56321 40371 56355
rect 40405 56352 40417 56355
rect 40862 56352 40868 56364
rect 40405 56324 40868 56352
rect 40405 56321 40417 56324
rect 40359 56315 40417 56321
rect 40862 56312 40868 56324
rect 40920 56312 40926 56364
rect 41046 56352 41052 56364
rect 41007 56324 41052 56352
rect 41046 56312 41052 56324
rect 41104 56312 41110 56364
rect 41233 56355 41291 56361
rect 41233 56321 41245 56355
rect 41279 56352 41291 56355
rect 41969 56355 42027 56361
rect 41969 56352 41981 56355
rect 41279 56324 41981 56352
rect 41279 56321 41291 56324
rect 41233 56315 41291 56321
rect 41969 56321 41981 56324
rect 42015 56321 42027 56355
rect 42150 56352 42156 56364
rect 42111 56324 42156 56352
rect 41969 56315 42027 56321
rect 42150 56312 42156 56324
rect 42208 56312 42214 56364
rect 42242 56312 42248 56364
rect 42300 56352 42306 56364
rect 42414 56355 42472 56361
rect 42300 56324 42345 56352
rect 42300 56312 42306 56324
rect 42414 56321 42426 56355
rect 42460 56321 42472 56355
rect 42414 56315 42472 56321
rect 40494 56284 40500 56296
rect 40455 56256 40500 56284
rect 40494 56244 40500 56256
rect 40552 56244 40558 56296
rect 40678 56244 40684 56296
rect 40736 56284 40742 56296
rect 41138 56284 41144 56296
rect 40736 56256 41144 56284
rect 40736 56244 40742 56256
rect 41138 56244 41144 56256
rect 41196 56244 41202 56296
rect 41414 56244 41420 56296
rect 41472 56284 41478 56296
rect 41509 56287 41567 56293
rect 41509 56284 41521 56287
rect 41472 56256 41521 56284
rect 41472 56244 41478 56256
rect 41509 56253 41521 56256
rect 41555 56253 41567 56287
rect 41509 56247 41567 56253
rect 41598 56244 41604 56296
rect 41656 56284 41662 56296
rect 42444 56284 42472 56315
rect 42518 56312 42524 56364
rect 42576 56352 42582 56364
rect 42576 56324 42621 56352
rect 42576 56312 42582 56324
rect 43070 56312 43076 56364
rect 43128 56352 43134 56364
rect 43257 56355 43315 56361
rect 43257 56352 43269 56355
rect 43128 56324 43269 56352
rect 43128 56312 43134 56324
rect 43257 56321 43269 56324
rect 43303 56321 43315 56355
rect 43530 56352 43536 56364
rect 43491 56324 43536 56352
rect 43257 56315 43315 56321
rect 43530 56312 43536 56324
rect 43588 56312 43594 56364
rect 43990 56312 43996 56364
rect 44048 56352 44054 56364
rect 44637 56355 44695 56361
rect 44637 56352 44649 56355
rect 44048 56324 44649 56352
rect 44048 56312 44054 56324
rect 44637 56321 44649 56324
rect 44683 56321 44695 56355
rect 44637 56315 44695 56321
rect 45462 56312 45468 56364
rect 45520 56352 45526 56364
rect 45556 56355 45614 56361
rect 45556 56352 45568 56355
rect 45520 56324 45568 56352
rect 45520 56312 45526 56324
rect 45556 56321 45568 56324
rect 45602 56321 45614 56355
rect 45556 56315 45614 56321
rect 45646 56312 45652 56364
rect 45704 56352 45710 56364
rect 45704 56324 45749 56352
rect 45704 56312 45710 56324
rect 46474 56312 46480 56364
rect 46532 56352 46538 56364
rect 47397 56355 47455 56361
rect 47397 56352 47409 56355
rect 46532 56324 47409 56352
rect 46532 56312 46538 56324
rect 47397 56321 47409 56324
rect 47443 56321 47455 56355
rect 47397 56315 47455 56321
rect 44542 56284 44548 56296
rect 41656 56256 42472 56284
rect 44503 56256 44548 56284
rect 41656 56244 41662 56256
rect 44542 56244 44548 56256
rect 44600 56244 44606 56296
rect 45094 56244 45100 56296
rect 45152 56284 45158 56296
rect 46753 56287 46811 56293
rect 46753 56284 46765 56287
rect 45152 56256 46765 56284
rect 45152 56244 45158 56256
rect 46753 56253 46765 56256
rect 46799 56253 46811 56287
rect 46753 56247 46811 56253
rect 43717 56219 43775 56225
rect 43717 56216 43729 56219
rect 38764 56188 40080 56216
rect 40144 56188 42472 56216
rect 26602 56148 26608 56160
rect 26160 56120 26608 56148
rect 26602 56108 26608 56120
rect 26660 56108 26666 56160
rect 27614 56108 27620 56160
rect 27672 56148 27678 56160
rect 29546 56148 29552 56160
rect 27672 56120 29552 56148
rect 27672 56108 27678 56120
rect 29546 56108 29552 56120
rect 29604 56108 29610 56160
rect 30650 56148 30656 56160
rect 30611 56120 30656 56148
rect 30650 56108 30656 56120
rect 30708 56108 30714 56160
rect 30926 56108 30932 56160
rect 30984 56148 30990 56160
rect 31846 56148 31852 56160
rect 30984 56120 31852 56148
rect 30984 56108 30990 56120
rect 31846 56108 31852 56120
rect 31904 56108 31910 56160
rect 33042 56108 33048 56160
rect 33100 56148 33106 56160
rect 33137 56151 33195 56157
rect 33137 56148 33149 56151
rect 33100 56120 33149 56148
rect 33100 56108 33106 56120
rect 33137 56117 33149 56120
rect 33183 56117 33195 56151
rect 33137 56111 33195 56117
rect 33318 56108 33324 56160
rect 33376 56148 33382 56160
rect 34517 56151 34575 56157
rect 34517 56148 34529 56151
rect 33376 56120 34529 56148
rect 33376 56108 33382 56120
rect 34517 56117 34529 56120
rect 34563 56148 34575 56151
rect 35710 56148 35716 56160
rect 34563 56120 35716 56148
rect 34563 56117 34575 56120
rect 34517 56111 34575 56117
rect 35710 56108 35716 56120
rect 35768 56108 35774 56160
rect 36630 56108 36636 56160
rect 36688 56148 36694 56160
rect 37645 56151 37703 56157
rect 37645 56148 37657 56151
rect 36688 56120 37657 56148
rect 36688 56108 36694 56120
rect 37645 56117 37657 56120
rect 37691 56117 37703 56151
rect 39850 56148 39856 56160
rect 39811 56120 39856 56148
rect 37645 56111 37703 56117
rect 39850 56108 39856 56120
rect 39908 56108 39914 56160
rect 40052 56148 40080 56188
rect 40678 56148 40684 56160
rect 40052 56120 40684 56148
rect 40678 56108 40684 56120
rect 40736 56108 40742 56160
rect 41414 56108 41420 56160
rect 41472 56148 41478 56160
rect 42444 56148 42472 56188
rect 42628 56188 43729 56216
rect 42628 56148 42656 56188
rect 43717 56185 43729 56188
rect 43763 56185 43775 56219
rect 43717 56179 43775 56185
rect 44634 56176 44640 56228
rect 44692 56216 44698 56228
rect 46109 56219 46167 56225
rect 44692 56188 45600 56216
rect 44692 56176 44698 56188
rect 41472 56120 41517 56148
rect 42444 56120 42656 56148
rect 41472 56108 41478 56120
rect 42886 56108 42892 56160
rect 42944 56148 42950 56160
rect 44361 56151 44419 56157
rect 44361 56148 44373 56151
rect 42944 56120 44373 56148
rect 42944 56108 42950 56120
rect 44361 56117 44373 56120
rect 44407 56117 44419 56151
rect 45462 56148 45468 56160
rect 45423 56120 45468 56148
rect 44361 56111 44419 56117
rect 45462 56108 45468 56120
rect 45520 56108 45526 56160
rect 45572 56148 45600 56188
rect 46109 56185 46121 56219
rect 46155 56185 46167 56219
rect 46109 56179 46167 56185
rect 46124 56148 46152 56179
rect 45572 56120 46152 56148
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 24765 55947 24823 55953
rect 24765 55913 24777 55947
rect 24811 55944 24823 55947
rect 25590 55944 25596 55956
rect 24811 55916 25596 55944
rect 24811 55913 24823 55916
rect 24765 55907 24823 55913
rect 25590 55904 25596 55916
rect 25648 55904 25654 55956
rect 26237 55947 26295 55953
rect 26237 55913 26249 55947
rect 26283 55944 26295 55947
rect 26326 55944 26332 55956
rect 26283 55916 26332 55944
rect 26283 55913 26295 55916
rect 26237 55907 26295 55913
rect 26326 55904 26332 55916
rect 26384 55904 26390 55956
rect 27709 55947 27767 55953
rect 27709 55913 27721 55947
rect 27755 55944 27767 55947
rect 30926 55944 30932 55956
rect 27755 55916 30932 55944
rect 27755 55913 27767 55916
rect 27709 55907 27767 55913
rect 30926 55904 30932 55916
rect 30984 55904 30990 55956
rect 33778 55904 33784 55956
rect 33836 55944 33842 55956
rect 35713 55947 35771 55953
rect 35713 55944 35725 55947
rect 33836 55916 35725 55944
rect 33836 55904 33842 55916
rect 35713 55913 35725 55916
rect 35759 55913 35771 55947
rect 35713 55907 35771 55913
rect 36722 55904 36728 55956
rect 36780 55944 36786 55956
rect 36817 55947 36875 55953
rect 36817 55944 36829 55947
rect 36780 55916 36829 55944
rect 36780 55904 36786 55916
rect 36817 55913 36829 55916
rect 36863 55913 36875 55947
rect 36817 55907 36875 55913
rect 37918 55904 37924 55956
rect 37976 55944 37982 55956
rect 38105 55947 38163 55953
rect 38105 55944 38117 55947
rect 37976 55916 38117 55944
rect 37976 55904 37982 55916
rect 38105 55913 38117 55916
rect 38151 55913 38163 55947
rect 38105 55907 38163 55913
rect 38286 55904 38292 55956
rect 38344 55944 38350 55956
rect 40221 55947 40279 55953
rect 40221 55944 40233 55947
rect 38344 55916 40233 55944
rect 38344 55904 38350 55916
rect 40221 55913 40233 55916
rect 40267 55913 40279 55947
rect 40221 55907 40279 55913
rect 40862 55904 40868 55956
rect 40920 55944 40926 55956
rect 41417 55947 41475 55953
rect 41417 55944 41429 55947
rect 40920 55916 41429 55944
rect 40920 55904 40926 55916
rect 41417 55913 41429 55916
rect 41463 55913 41475 55947
rect 41417 55907 41475 55913
rect 42337 55947 42395 55953
rect 42337 55913 42349 55947
rect 42383 55944 42395 55947
rect 42518 55944 42524 55956
rect 42383 55916 42524 55944
rect 42383 55913 42395 55916
rect 42337 55907 42395 55913
rect 42518 55904 42524 55916
rect 42576 55904 42582 55956
rect 42705 55947 42763 55953
rect 42705 55913 42717 55947
rect 42751 55944 42763 55947
rect 43162 55944 43168 55956
rect 42751 55916 43168 55944
rect 42751 55913 42763 55916
rect 42705 55907 42763 55913
rect 43162 55904 43168 55916
rect 43220 55904 43226 55956
rect 44542 55904 44548 55956
rect 44600 55944 44606 55956
rect 44637 55947 44695 55953
rect 44637 55944 44649 55947
rect 44600 55916 44649 55944
rect 44600 55904 44606 55916
rect 44637 55913 44649 55916
rect 44683 55913 44695 55947
rect 46750 55944 46756 55956
rect 44637 55907 44695 55913
rect 44836 55916 46756 55944
rect 26878 55876 26884 55888
rect 26791 55848 26884 55876
rect 26878 55836 26884 55848
rect 26936 55876 26942 55888
rect 31481 55879 31539 55885
rect 31481 55876 31493 55879
rect 26936 55848 31493 55876
rect 26936 55836 26942 55848
rect 31481 55845 31493 55848
rect 31527 55845 31539 55879
rect 31481 55839 31539 55845
rect 34701 55879 34759 55885
rect 34701 55845 34713 55879
rect 34747 55845 34759 55879
rect 34701 55839 34759 55845
rect 23201 55811 23259 55817
rect 23201 55777 23213 55811
rect 23247 55808 23259 55811
rect 23661 55811 23719 55817
rect 23661 55808 23673 55811
rect 23247 55780 23673 55808
rect 23247 55777 23259 55780
rect 23201 55771 23259 55777
rect 23661 55777 23673 55780
rect 23707 55808 23719 55811
rect 24762 55808 24768 55820
rect 23707 55780 24768 55808
rect 23707 55777 23719 55780
rect 23661 55771 23719 55777
rect 24762 55768 24768 55780
rect 24820 55768 24826 55820
rect 23750 55700 23756 55752
rect 23808 55740 23814 55752
rect 23845 55743 23903 55749
rect 23845 55740 23857 55743
rect 23808 55712 23857 55740
rect 23808 55700 23814 55712
rect 23845 55709 23857 55712
rect 23891 55709 23903 55743
rect 23845 55703 23903 55709
rect 24581 55743 24639 55749
rect 24581 55709 24593 55743
rect 24627 55740 24639 55743
rect 25225 55743 25283 55749
rect 25225 55740 25237 55743
rect 24627 55712 25237 55740
rect 24627 55709 24639 55712
rect 24581 55703 24639 55709
rect 25225 55709 25237 55712
rect 25271 55709 25283 55743
rect 25225 55703 25283 55709
rect 25406 55700 25412 55752
rect 25464 55740 25470 55752
rect 26896 55749 26924 55836
rect 28258 55808 28264 55820
rect 26988 55780 28264 55808
rect 26988 55752 27016 55780
rect 28258 55768 28264 55780
rect 28316 55768 28322 55820
rect 28442 55808 28448 55820
rect 28403 55780 28448 55808
rect 28442 55768 28448 55780
rect 28500 55768 28506 55820
rect 28534 55768 28540 55820
rect 28592 55808 28598 55820
rect 28721 55811 28779 55817
rect 28721 55808 28733 55811
rect 28592 55780 28733 55808
rect 28592 55768 28598 55780
rect 28721 55777 28733 55780
rect 28767 55777 28779 55811
rect 28721 55771 28779 55777
rect 28905 55811 28963 55817
rect 28905 55777 28917 55811
rect 28951 55808 28963 55811
rect 29362 55808 29368 55820
rect 28951 55780 29368 55808
rect 28951 55777 28963 55780
rect 28905 55771 28963 55777
rect 29362 55768 29368 55780
rect 29420 55768 29426 55820
rect 29914 55808 29920 55820
rect 29656 55780 29920 55808
rect 25593 55743 25651 55749
rect 25464 55712 25557 55740
rect 25464 55700 25470 55712
rect 25593 55709 25605 55743
rect 25639 55709 25651 55743
rect 25593 55703 25651 55709
rect 26053 55743 26111 55749
rect 26053 55709 26065 55743
rect 26099 55740 26111 55743
rect 26697 55743 26755 55749
rect 26697 55740 26709 55743
rect 26099 55712 26709 55740
rect 26099 55709 26111 55712
rect 26053 55703 26111 55709
rect 26697 55709 26709 55712
rect 26743 55709 26755 55743
rect 26697 55703 26755 55709
rect 26881 55743 26939 55749
rect 26881 55709 26893 55743
rect 26927 55709 26939 55743
rect 26881 55703 26939 55709
rect 24026 55604 24032 55616
rect 23987 55576 24032 55604
rect 24026 55564 24032 55576
rect 24084 55564 24090 55616
rect 25424 55604 25452 55700
rect 25608 55672 25636 55703
rect 26970 55700 26976 55752
rect 27028 55740 27034 55752
rect 27525 55743 27583 55749
rect 27028 55712 27073 55740
rect 27028 55700 27034 55712
rect 27525 55709 27537 55743
rect 27571 55709 27583 55743
rect 28626 55740 28632 55752
rect 28587 55712 28632 55740
rect 27525 55703 27583 55709
rect 26988 55672 27016 55700
rect 25608 55644 27016 55672
rect 27540 55672 27568 55703
rect 28626 55700 28632 55712
rect 28684 55700 28690 55752
rect 28810 55740 28816 55752
rect 28771 55712 28816 55740
rect 28810 55700 28816 55712
rect 28868 55700 28874 55752
rect 29656 55749 29684 55780
rect 29914 55768 29920 55780
rect 29972 55808 29978 55820
rect 34716 55808 34744 55839
rect 35526 55836 35532 55888
rect 35584 55876 35590 55888
rect 37369 55879 37427 55885
rect 37369 55876 37381 55879
rect 35584 55848 37381 55876
rect 35584 55836 35590 55848
rect 37369 55845 37381 55848
rect 37415 55845 37427 55879
rect 37369 55839 37427 55845
rect 34974 55808 34980 55820
rect 29972 55780 34744 55808
rect 34935 55780 34980 55808
rect 29972 55768 29978 55780
rect 34974 55768 34980 55780
rect 35032 55768 35038 55820
rect 36630 55808 36636 55820
rect 36591 55780 36636 55808
rect 36630 55768 36636 55780
rect 36688 55768 36694 55820
rect 38304 55808 38332 55904
rect 38378 55836 38384 55888
rect 38436 55836 38442 55888
rect 38562 55876 38568 55888
rect 38488 55848 38568 55876
rect 37568 55780 38332 55808
rect 29641 55743 29699 55749
rect 29641 55709 29653 55743
rect 29687 55709 29699 55743
rect 29641 55703 29699 55709
rect 29730 55700 29736 55752
rect 29788 55740 29794 55752
rect 29825 55743 29883 55749
rect 29825 55740 29837 55743
rect 29788 55712 29837 55740
rect 29788 55700 29794 55712
rect 29825 55709 29837 55712
rect 29871 55740 29883 55743
rect 30098 55740 30104 55752
rect 29871 55712 30104 55740
rect 29871 55709 29883 55712
rect 29825 55703 29883 55709
rect 30098 55700 30104 55712
rect 30156 55700 30162 55752
rect 30834 55740 30840 55752
rect 30795 55712 30840 55740
rect 30834 55700 30840 55712
rect 30892 55700 30898 55752
rect 31294 55740 31300 55752
rect 31255 55712 31300 55740
rect 31294 55700 31300 55712
rect 31352 55700 31358 55752
rect 32125 55743 32183 55749
rect 32125 55709 32137 55743
rect 32171 55709 32183 55743
rect 32398 55740 32404 55752
rect 32311 55712 32404 55740
rect 32125 55703 32183 55709
rect 27890 55672 27896 55684
rect 27540 55644 27896 55672
rect 27890 55632 27896 55644
rect 27948 55672 27954 55684
rect 28994 55672 29000 55684
rect 27948 55644 29000 55672
rect 27948 55632 27954 55644
rect 28994 55632 29000 55644
rect 29052 55632 29058 55684
rect 30742 55632 30748 55684
rect 30800 55672 30806 55684
rect 30975 55675 31033 55681
rect 30975 55672 30987 55675
rect 30800 55644 30987 55672
rect 30800 55632 30806 55644
rect 30975 55641 30987 55644
rect 31021 55641 31033 55675
rect 31110 55672 31116 55684
rect 31071 55644 31116 55672
rect 30975 55635 31033 55641
rect 31110 55632 31116 55644
rect 31168 55632 31174 55684
rect 31205 55675 31263 55681
rect 31205 55641 31217 55675
rect 31251 55672 31263 55675
rect 31941 55675 31999 55681
rect 31941 55672 31953 55675
rect 31251 55644 31953 55672
rect 31251 55641 31263 55644
rect 31205 55635 31263 55641
rect 31941 55641 31953 55644
rect 31987 55641 31999 55675
rect 32140 55672 32168 55703
rect 32398 55700 32404 55712
rect 32456 55740 32462 55752
rect 32674 55740 32680 55752
rect 32456 55712 32680 55740
rect 32456 55700 32462 55712
rect 32674 55700 32680 55712
rect 32732 55700 32738 55752
rect 33042 55740 33048 55752
rect 33003 55712 33048 55740
rect 33042 55700 33048 55712
rect 33100 55700 33106 55752
rect 33226 55740 33232 55752
rect 33187 55712 33232 55740
rect 33226 55700 33232 55712
rect 33284 55700 33290 55752
rect 33321 55743 33379 55749
rect 33321 55709 33333 55743
rect 33367 55740 33379 55743
rect 33686 55740 33692 55752
rect 33367 55712 33692 55740
rect 33367 55709 33379 55712
rect 33321 55703 33379 55709
rect 33686 55700 33692 55712
rect 33744 55700 33750 55752
rect 34054 55700 34060 55752
rect 34112 55740 34118 55752
rect 34790 55740 34796 55752
rect 34112 55712 34796 55740
rect 34112 55700 34118 55712
rect 34790 55700 34796 55712
rect 34848 55700 34854 55752
rect 35069 55743 35127 55749
rect 35069 55709 35081 55743
rect 35115 55740 35127 55743
rect 36078 55740 36084 55752
rect 35115 55712 36084 55740
rect 35115 55709 35127 55712
rect 35069 55703 35127 55709
rect 32858 55672 32864 55684
rect 32140 55644 32444 55672
rect 32819 55644 32864 55672
rect 31941 55635 31999 55641
rect 29270 55604 29276 55616
rect 25424 55576 29276 55604
rect 29270 55564 29276 55576
rect 29328 55564 29334 55616
rect 29454 55604 29460 55616
rect 29415 55576 29460 55604
rect 29454 55564 29460 55576
rect 29512 55564 29518 55616
rect 30377 55607 30435 55613
rect 30377 55573 30389 55607
rect 30423 55604 30435 55607
rect 30650 55604 30656 55616
rect 30423 55576 30656 55604
rect 30423 55573 30435 55576
rect 30377 55567 30435 55573
rect 30650 55564 30656 55576
rect 30708 55604 30714 55616
rect 31128 55604 31156 55632
rect 32306 55604 32312 55616
rect 30708 55576 31156 55604
rect 32267 55576 32312 55604
rect 30708 55564 30714 55576
rect 32306 55564 32312 55576
rect 32364 55564 32370 55616
rect 32416 55604 32444 55644
rect 32858 55632 32864 55644
rect 32916 55632 32922 55684
rect 34330 55632 34336 55684
rect 34388 55672 34394 55684
rect 35084 55672 35112 55703
rect 36078 55700 36084 55712
rect 36136 55700 36142 55752
rect 36538 55740 36544 55752
rect 36499 55712 36544 55740
rect 36538 55700 36544 55712
rect 36596 55700 36602 55752
rect 37568 55749 37596 55780
rect 37553 55743 37611 55749
rect 37553 55709 37565 55743
rect 37599 55709 37611 55743
rect 37553 55703 37611 55709
rect 37645 55743 37703 55749
rect 37645 55709 37657 55743
rect 37691 55740 37703 55743
rect 37918 55740 37924 55752
rect 37691 55712 37924 55740
rect 37691 55709 37703 55712
rect 37645 55703 37703 55709
rect 37918 55700 37924 55712
rect 37976 55700 37982 55752
rect 38286 55740 38292 55752
rect 38247 55712 38292 55740
rect 38286 55700 38292 55712
rect 38344 55700 38350 55752
rect 38396 55749 38424 55836
rect 38381 55743 38439 55749
rect 38381 55709 38393 55743
rect 38427 55709 38439 55743
rect 38488 55740 38516 55848
rect 38562 55836 38568 55848
rect 38620 55836 38626 55888
rect 38930 55836 38936 55888
rect 38988 55876 38994 55888
rect 40402 55876 40408 55888
rect 38988 55848 40408 55876
rect 38988 55836 38994 55848
rect 40402 55836 40408 55848
rect 40460 55876 40466 55888
rect 40770 55876 40776 55888
rect 40460 55848 40776 55876
rect 40460 55836 40466 55848
rect 40770 55836 40776 55848
rect 40828 55836 40834 55888
rect 40954 55836 40960 55888
rect 41012 55876 41018 55888
rect 41690 55876 41696 55888
rect 41012 55848 41696 55876
rect 41012 55836 41018 55848
rect 41690 55836 41696 55848
rect 41748 55836 41754 55888
rect 42242 55836 42248 55888
rect 42300 55876 42306 55888
rect 42794 55876 42800 55888
rect 42300 55848 42800 55876
rect 42300 55836 42306 55848
rect 42794 55836 42800 55848
rect 42852 55836 42858 55888
rect 44177 55879 44235 55885
rect 44177 55876 44189 55879
rect 43364 55848 44189 55876
rect 40586 55768 40592 55820
rect 40644 55808 40650 55820
rect 43257 55811 43315 55817
rect 43257 55808 43269 55811
rect 40644 55780 43269 55808
rect 40644 55768 40650 55780
rect 43257 55777 43269 55780
rect 43303 55777 43315 55811
rect 43257 55771 43315 55777
rect 38565 55743 38623 55749
rect 38565 55740 38577 55743
rect 38488 55712 38577 55740
rect 38381 55703 38439 55709
rect 38565 55709 38577 55712
rect 38611 55709 38623 55743
rect 38565 55703 38623 55709
rect 38654 55700 38660 55752
rect 38712 55740 38718 55752
rect 39298 55740 39304 55752
rect 38712 55712 38757 55740
rect 39259 55712 39304 55740
rect 38712 55700 38718 55712
rect 39298 55700 39304 55712
rect 39356 55700 39362 55752
rect 39482 55740 39488 55752
rect 39443 55712 39488 55740
rect 39482 55700 39488 55712
rect 39540 55700 39546 55752
rect 39942 55700 39948 55752
rect 40000 55740 40006 55752
rect 40000 55712 40724 55740
rect 40000 55700 40006 55712
rect 34388 55644 35112 55672
rect 37369 55675 37427 55681
rect 34388 55632 34394 55644
rect 37369 55641 37381 55675
rect 37415 55641 37427 55675
rect 39114 55672 39120 55684
rect 39075 55644 39120 55672
rect 37369 55635 37427 55641
rect 35158 55604 35164 55616
rect 32416 55576 35164 55604
rect 35158 55564 35164 55576
rect 35216 55564 35222 55616
rect 37384 55604 37412 55635
rect 39114 55632 39120 55644
rect 39172 55632 39178 55684
rect 40402 55672 40408 55684
rect 40363 55644 40408 55672
rect 40402 55632 40408 55644
rect 40460 55632 40466 55684
rect 40586 55672 40592 55684
rect 40547 55644 40592 55672
rect 40586 55632 40592 55644
rect 40644 55632 40650 55684
rect 40696 55672 40724 55712
rect 40862 55700 40868 55752
rect 40920 55740 40926 55752
rect 41049 55743 41107 55749
rect 41049 55740 41061 55743
rect 40920 55712 41061 55740
rect 40920 55700 40926 55712
rect 41049 55709 41061 55712
rect 41095 55709 41107 55743
rect 41049 55703 41107 55709
rect 42521 55743 42579 55749
rect 42521 55709 42533 55743
rect 42567 55740 42579 55743
rect 42610 55740 42616 55752
rect 42567 55712 42616 55740
rect 42567 55709 42579 55712
rect 42521 55703 42579 55709
rect 42610 55700 42616 55712
rect 42668 55700 42674 55752
rect 42794 55740 42800 55752
rect 42755 55712 42800 55740
rect 42794 55700 42800 55712
rect 42852 55700 42858 55752
rect 41233 55675 41291 55681
rect 41233 55672 41245 55675
rect 40696 55644 41245 55672
rect 41233 55641 41245 55644
rect 41279 55641 41291 55675
rect 41233 55635 41291 55641
rect 41322 55632 41328 55684
rect 41380 55672 41386 55684
rect 43364 55672 43392 55848
rect 44177 55845 44189 55848
rect 44223 55845 44235 55879
rect 44177 55839 44235 55845
rect 44266 55836 44272 55888
rect 44324 55876 44330 55888
rect 44836 55876 44864 55916
rect 46750 55904 46756 55916
rect 46808 55904 46814 55956
rect 46934 55904 46940 55956
rect 46992 55944 46998 55956
rect 47305 55947 47363 55953
rect 47305 55944 47317 55947
rect 46992 55916 47317 55944
rect 46992 55904 46998 55916
rect 47305 55913 47317 55916
rect 47351 55913 47363 55947
rect 47305 55907 47363 55913
rect 45002 55876 45008 55888
rect 44324 55848 44864 55876
rect 44963 55848 45008 55876
rect 44324 55836 44330 55848
rect 45002 55836 45008 55848
rect 45060 55836 45066 55888
rect 45646 55836 45652 55888
rect 45704 55876 45710 55888
rect 46293 55879 46351 55885
rect 46293 55876 46305 55879
rect 45704 55848 46305 55876
rect 45704 55836 45710 55848
rect 46293 55845 46305 55848
rect 46339 55876 46351 55879
rect 55398 55876 55404 55888
rect 46339 55848 55404 55876
rect 46339 55845 46351 55848
rect 46293 55839 46351 55845
rect 55398 55836 55404 55848
rect 55456 55836 55462 55888
rect 43530 55768 43536 55820
rect 43588 55808 43594 55820
rect 47486 55808 47492 55820
rect 43588 55780 47492 55808
rect 43588 55768 43594 55780
rect 43901 55743 43959 55749
rect 43901 55709 43913 55743
rect 43947 55709 43959 55743
rect 43901 55703 43959 55709
rect 41380 55644 43392 55672
rect 43916 55672 43944 55703
rect 43990 55700 43996 55752
rect 44048 55740 44054 55752
rect 44177 55743 44235 55749
rect 44048 55712 44093 55740
rect 44048 55700 44054 55712
rect 44177 55709 44189 55743
rect 44223 55740 44235 55743
rect 44542 55740 44548 55752
rect 44223 55712 44548 55740
rect 44223 55709 44235 55712
rect 44177 55703 44235 55709
rect 44542 55700 44548 55712
rect 44600 55700 44606 55752
rect 44836 55749 44864 55780
rect 47486 55768 47492 55780
rect 47544 55768 47550 55820
rect 44821 55743 44879 55749
rect 44821 55709 44833 55743
rect 44867 55709 44879 55743
rect 44821 55703 44879 55709
rect 44910 55700 44916 55752
rect 44968 55740 44974 55752
rect 45097 55743 45155 55749
rect 44968 55712 45013 55740
rect 44968 55700 44974 55712
rect 45097 55709 45109 55743
rect 45143 55740 45155 55743
rect 45462 55740 45468 55752
rect 45143 55712 45468 55740
rect 45143 55709 45155 55712
rect 45097 55703 45155 55709
rect 44726 55672 44732 55684
rect 43916 55644 44732 55672
rect 41380 55632 41386 55644
rect 44726 55632 44732 55644
rect 44784 55672 44790 55684
rect 45112 55672 45140 55703
rect 45462 55700 45468 55712
rect 45520 55700 45526 55752
rect 44784 55644 45140 55672
rect 44784 55632 44790 55644
rect 38102 55604 38108 55616
rect 37384 55576 38108 55604
rect 38102 55564 38108 55576
rect 38160 55604 38166 55616
rect 40678 55604 40684 55616
rect 38160 55576 40684 55604
rect 38160 55564 38166 55576
rect 40678 55564 40684 55576
rect 40736 55564 40742 55616
rect 40770 55564 40776 55616
rect 40828 55604 40834 55616
rect 42886 55604 42892 55616
rect 40828 55576 42892 55604
rect 40828 55564 40834 55576
rect 42886 55564 42892 55576
rect 42944 55564 42950 55616
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 23382 55360 23388 55412
rect 23440 55400 23446 55412
rect 23845 55403 23903 55409
rect 23845 55400 23857 55403
rect 23440 55372 23857 55400
rect 23440 55360 23446 55372
rect 23845 55369 23857 55372
rect 23891 55369 23903 55403
rect 23845 55363 23903 55369
rect 25501 55403 25559 55409
rect 25501 55369 25513 55403
rect 25547 55400 25559 55403
rect 25774 55400 25780 55412
rect 25547 55372 25780 55400
rect 25547 55369 25559 55372
rect 25501 55363 25559 55369
rect 25774 55360 25780 55372
rect 25832 55360 25838 55412
rect 26234 55400 26240 55412
rect 26195 55372 26240 55400
rect 26234 55360 26240 55372
rect 26292 55360 26298 55412
rect 28350 55360 28356 55412
rect 28408 55400 28414 55412
rect 28810 55400 28816 55412
rect 28408 55372 28816 55400
rect 28408 55360 28414 55372
rect 28810 55360 28816 55372
rect 28868 55400 28874 55412
rect 30742 55400 30748 55412
rect 28868 55372 29684 55400
rect 30703 55372 30748 55400
rect 28868 55360 28874 55372
rect 28997 55335 29055 55341
rect 28997 55301 29009 55335
rect 29043 55332 29055 55335
rect 29454 55332 29460 55344
rect 29043 55304 29460 55332
rect 29043 55301 29055 55304
rect 28997 55295 29055 55301
rect 29454 55292 29460 55304
rect 29512 55292 29518 55344
rect 24026 55264 24032 55276
rect 23987 55236 24032 55264
rect 24026 55224 24032 55236
rect 24084 55224 24090 55276
rect 25682 55264 25688 55276
rect 25643 55236 25688 55264
rect 25682 55224 25688 55236
rect 25740 55224 25746 55276
rect 26418 55264 26424 55276
rect 26379 55236 26424 55264
rect 26418 55224 26424 55236
rect 26476 55224 26482 55276
rect 26602 55224 26608 55276
rect 26660 55264 26666 55276
rect 26881 55267 26939 55273
rect 26881 55264 26893 55267
rect 26660 55236 26893 55264
rect 26660 55224 26666 55236
rect 26881 55233 26893 55236
rect 26927 55233 26939 55267
rect 26881 55227 26939 55233
rect 26973 55267 27031 55273
rect 26973 55233 26985 55267
rect 27019 55264 27031 55267
rect 27522 55264 27528 55276
rect 27019 55236 27528 55264
rect 27019 55233 27031 55236
rect 26973 55227 27031 55233
rect 27522 55224 27528 55236
rect 27580 55224 27586 55276
rect 27706 55264 27712 55276
rect 27667 55236 27712 55264
rect 27706 55224 27712 55236
rect 27764 55224 27770 55276
rect 27801 55267 27859 55273
rect 27801 55233 27813 55267
rect 27847 55264 27859 55267
rect 28442 55264 28448 55276
rect 27847 55236 28448 55264
rect 27847 55233 27859 55236
rect 27801 55227 27859 55233
rect 28442 55224 28448 55236
rect 28500 55224 28506 55276
rect 29549 55267 29607 55273
rect 29549 55264 29561 55267
rect 28644 55236 29561 55264
rect 28534 55156 28540 55208
rect 28592 55196 28598 55208
rect 28644 55196 28672 55236
rect 29549 55233 29561 55236
rect 29595 55233 29607 55267
rect 29656 55264 29684 55372
rect 30742 55360 30748 55372
rect 30800 55360 30806 55412
rect 31294 55360 31300 55412
rect 31352 55400 31358 55412
rect 33045 55403 33103 55409
rect 33045 55400 33057 55403
rect 31352 55372 33057 55400
rect 31352 55360 31358 55372
rect 33045 55369 33057 55372
rect 33091 55369 33103 55403
rect 34418 55403 34476 55409
rect 34418 55400 34430 55403
rect 33045 55363 33103 55369
rect 33152 55372 34430 55400
rect 29730 55292 29736 55344
rect 29788 55332 29794 55344
rect 29914 55332 29920 55344
rect 29788 55304 29833 55332
rect 29875 55304 29920 55332
rect 29788 55292 29794 55304
rect 29914 55292 29920 55304
rect 29972 55292 29978 55344
rect 33152 55332 33180 55372
rect 34418 55369 34430 55372
rect 34464 55369 34476 55403
rect 34974 55400 34980 55412
rect 34418 55363 34476 55369
rect 34532 55372 34980 55400
rect 33594 55332 33600 55344
rect 30024 55304 33180 55332
rect 33555 55304 33600 55332
rect 30024 55264 30052 55304
rect 33594 55292 33600 55304
rect 33652 55292 33658 55344
rect 34330 55332 34336 55344
rect 34291 55304 34336 55332
rect 34330 55292 34336 55304
rect 34388 55292 34394 55344
rect 34532 55341 34560 55372
rect 34974 55360 34980 55372
rect 35032 55360 35038 55412
rect 35158 55360 35164 55412
rect 35216 55400 35222 55412
rect 35434 55400 35440 55412
rect 35216 55372 35440 55400
rect 35216 55360 35222 55372
rect 35434 55360 35440 55372
rect 35492 55360 35498 55412
rect 36538 55360 36544 55412
rect 36596 55400 36602 55412
rect 38105 55403 38163 55409
rect 38105 55400 38117 55403
rect 36596 55372 38117 55400
rect 36596 55360 36602 55372
rect 38105 55369 38117 55372
rect 38151 55369 38163 55403
rect 38105 55363 38163 55369
rect 38378 55360 38384 55412
rect 38436 55400 38442 55412
rect 38473 55403 38531 55409
rect 38473 55400 38485 55403
rect 38436 55372 38485 55400
rect 38436 55360 38442 55372
rect 38473 55369 38485 55372
rect 38519 55400 38531 55403
rect 39114 55400 39120 55412
rect 38519 55372 39120 55400
rect 38519 55369 38531 55372
rect 38473 55363 38531 55369
rect 39114 55360 39120 55372
rect 39172 55360 39178 55412
rect 40030 55403 40088 55409
rect 40030 55369 40042 55403
rect 40076 55400 40088 55403
rect 40494 55400 40500 55412
rect 40076 55372 40500 55400
rect 40076 55369 40088 55372
rect 40030 55363 40088 55369
rect 40494 55360 40500 55372
rect 40552 55360 40558 55412
rect 40678 55360 40684 55412
rect 40736 55400 40742 55412
rect 41230 55400 41236 55412
rect 40736 55372 41236 55400
rect 40736 55360 40742 55372
rect 41230 55360 41236 55372
rect 41288 55360 41294 55412
rect 42426 55360 42432 55412
rect 42484 55400 42490 55412
rect 42484 55372 44036 55400
rect 42484 55360 42490 55372
rect 34517 55335 34575 55341
rect 34517 55301 34529 55335
rect 34563 55301 34575 55335
rect 34517 55295 34575 55301
rect 34606 55292 34612 55344
rect 34664 55332 34670 55344
rect 34664 55304 35388 55332
rect 34664 55292 34670 55304
rect 30374 55264 30380 55276
rect 29656 55236 30052 55264
rect 30335 55236 30380 55264
rect 29549 55227 29607 55233
rect 30374 55224 30380 55236
rect 30432 55224 30438 55276
rect 30558 55264 30564 55276
rect 30519 55236 30564 55264
rect 30558 55224 30564 55236
rect 30616 55224 30622 55276
rect 31570 55224 31576 55276
rect 31628 55264 31634 55276
rect 31757 55267 31815 55273
rect 31757 55264 31769 55267
rect 31628 55236 31769 55264
rect 31628 55224 31634 55236
rect 31757 55233 31769 55236
rect 31803 55233 31815 55267
rect 32674 55264 32680 55276
rect 32635 55236 32680 55264
rect 31757 55227 31815 55233
rect 32674 55224 32680 55236
rect 32732 55224 32738 55276
rect 32861 55267 32919 55273
rect 32861 55233 32873 55267
rect 32907 55264 32919 55267
rect 33318 55264 33324 55276
rect 32907 55236 33324 55264
rect 32907 55233 32919 55236
rect 32861 55227 32919 55233
rect 28592 55168 28672 55196
rect 28592 55156 28598 55168
rect 28644 55137 28672 55168
rect 32306 55156 32312 55208
rect 32364 55196 32370 55208
rect 32876 55196 32904 55227
rect 33318 55224 33324 55236
rect 33376 55224 33382 55276
rect 33686 55264 33692 55276
rect 33647 55236 33692 55264
rect 33686 55224 33692 55236
rect 33744 55224 33750 55276
rect 34241 55267 34299 55273
rect 34241 55233 34253 55267
rect 34287 55233 34299 55267
rect 35158 55264 35164 55276
rect 35119 55236 35164 55264
rect 34241 55227 34299 55233
rect 32364 55168 32904 55196
rect 34256 55196 34284 55227
rect 35158 55224 35164 55236
rect 35216 55224 35222 55276
rect 35360 55273 35388 55304
rect 35618 55292 35624 55344
rect 35676 55332 35682 55344
rect 38654 55332 38660 55344
rect 35676 55304 37320 55332
rect 35676 55292 35682 55304
rect 35345 55267 35403 55273
rect 35345 55233 35357 55267
rect 35391 55233 35403 55267
rect 35345 55227 35403 55233
rect 35437 55267 35495 55273
rect 35437 55233 35449 55267
rect 35483 55233 35495 55267
rect 35437 55227 35495 55233
rect 34422 55196 34428 55208
rect 34256 55168 34428 55196
rect 32364 55156 32370 55168
rect 34422 55156 34428 55168
rect 34480 55196 34486 55208
rect 35452 55196 35480 55227
rect 35526 55224 35532 55276
rect 35584 55264 35590 55276
rect 35710 55264 35716 55276
rect 35584 55236 35716 55264
rect 35584 55224 35590 55236
rect 35710 55224 35716 55236
rect 35768 55264 35774 55276
rect 36264 55267 36322 55273
rect 36264 55264 36276 55267
rect 35768 55236 36276 55264
rect 35768 55224 35774 55236
rect 36264 55233 36276 55236
rect 36310 55233 36322 55267
rect 36264 55227 36322 55233
rect 36357 55267 36415 55273
rect 36357 55233 36369 55267
rect 36403 55264 36415 55267
rect 36446 55264 36452 55276
rect 36403 55236 36452 55264
rect 36403 55233 36415 55236
rect 36357 55227 36415 55233
rect 35989 55199 36047 55205
rect 35989 55196 36001 55199
rect 34480 55168 36001 55196
rect 34480 55156 34486 55168
rect 35989 55165 36001 55168
rect 36035 55165 36047 55199
rect 35989 55159 36047 55165
rect 28629 55131 28687 55137
rect 28629 55097 28641 55131
rect 28675 55097 28687 55131
rect 28629 55091 28687 55097
rect 34882 55088 34888 55140
rect 34940 55128 34946 55140
rect 35253 55131 35311 55137
rect 35253 55128 35265 55131
rect 34940 55100 35265 55128
rect 34940 55088 34946 55100
rect 35253 55097 35265 55100
rect 35299 55128 35311 55131
rect 35710 55128 35716 55140
rect 35299 55100 35716 55128
rect 35299 55097 35311 55100
rect 35253 55091 35311 55097
rect 35710 55088 35716 55100
rect 35768 55088 35774 55140
rect 36279 55128 36307 55227
rect 36446 55224 36452 55236
rect 36504 55224 36510 55276
rect 37292 55205 37320 55304
rect 38304 55304 38660 55332
rect 38304 55273 38332 55304
rect 38654 55292 38660 55304
rect 38712 55332 38718 55344
rect 39025 55335 39083 55341
rect 39025 55332 39037 55335
rect 38712 55304 39037 55332
rect 38712 55292 38718 55304
rect 39025 55301 39037 55304
rect 39071 55301 39083 55335
rect 39942 55332 39948 55344
rect 39025 55295 39083 55301
rect 39132 55304 39804 55332
rect 39903 55304 39948 55332
rect 38289 55267 38347 55273
rect 38289 55233 38301 55267
rect 38335 55233 38347 55267
rect 38289 55227 38347 55233
rect 38378 55224 38384 55276
rect 38436 55264 38442 55276
rect 38565 55267 38623 55273
rect 38565 55264 38577 55267
rect 38436 55236 38577 55264
rect 38436 55224 38442 55236
rect 38565 55233 38577 55236
rect 38611 55264 38623 55267
rect 39132 55264 39160 55304
rect 38611 55236 39160 55264
rect 39209 55267 39267 55273
rect 38611 55233 38623 55236
rect 38565 55227 38623 55233
rect 39209 55233 39221 55267
rect 39255 55264 39267 55267
rect 39482 55264 39488 55276
rect 39255 55236 39488 55264
rect 39255 55233 39267 55236
rect 39209 55227 39267 55233
rect 39482 55224 39488 55236
rect 39540 55224 39546 55276
rect 39776 55264 39804 55304
rect 39942 55292 39948 55304
rect 40000 55292 40006 55344
rect 40129 55335 40187 55341
rect 40129 55301 40141 55335
rect 40175 55332 40187 55335
rect 40218 55332 40224 55344
rect 40175 55304 40224 55332
rect 40175 55301 40187 55304
rect 40129 55295 40187 55301
rect 40218 55292 40224 55304
rect 40276 55292 40282 55344
rect 44008 55341 44036 55372
rect 44082 55360 44088 55412
rect 44140 55400 44146 55412
rect 44453 55403 44511 55409
rect 44453 55400 44465 55403
rect 44140 55372 44465 55400
rect 44140 55360 44146 55372
rect 44453 55369 44465 55372
rect 44499 55369 44511 55403
rect 44453 55363 44511 55369
rect 45097 55403 45155 55409
rect 45097 55369 45109 55403
rect 45143 55400 45155 55403
rect 45186 55400 45192 55412
rect 45143 55372 45192 55400
rect 45143 55369 45155 55372
rect 45097 55363 45155 55369
rect 45186 55360 45192 55372
rect 45244 55360 45250 55412
rect 45554 55400 45560 55412
rect 45515 55372 45560 55400
rect 45554 55360 45560 55372
rect 45612 55360 45618 55412
rect 43993 55335 44051 55341
rect 43993 55301 44005 55335
rect 44039 55332 44051 55335
rect 45646 55332 45652 55344
rect 44039 55304 45652 55332
rect 44039 55301 44051 55304
rect 43993 55295 44051 55301
rect 45646 55292 45652 55304
rect 45704 55292 45710 55344
rect 39850 55264 39856 55276
rect 39763 55236 39856 55264
rect 39850 55224 39856 55236
rect 39908 55224 39914 55276
rect 40681 55267 40739 55273
rect 40681 55233 40693 55267
rect 40727 55233 40739 55267
rect 40681 55227 40739 55233
rect 37277 55199 37335 55205
rect 37277 55165 37289 55199
rect 37323 55165 37335 55199
rect 37277 55159 37335 55165
rect 39298 55156 39304 55208
rect 39356 55196 39362 55208
rect 39393 55199 39451 55205
rect 39393 55196 39405 55199
rect 39356 55168 39405 55196
rect 39356 55156 39362 55168
rect 39393 55165 39405 55168
rect 39439 55165 39451 55199
rect 39393 55159 39451 55165
rect 40696 55128 40724 55227
rect 41966 55224 41972 55276
rect 42024 55264 42030 55276
rect 42061 55267 42119 55273
rect 42061 55264 42073 55267
rect 42024 55236 42073 55264
rect 42024 55224 42030 55236
rect 42061 55233 42073 55236
rect 42107 55233 42119 55267
rect 42061 55227 42119 55233
rect 42334 55224 42340 55276
rect 42392 55264 42398 55276
rect 42392 55236 43300 55264
rect 42392 55224 42398 55236
rect 41138 55156 41144 55208
rect 41196 55156 41202 55208
rect 41874 55156 41880 55208
rect 41932 55196 41938 55208
rect 43272 55205 43300 55236
rect 42521 55199 42579 55205
rect 42521 55196 42533 55199
rect 41932 55168 42533 55196
rect 41932 55156 41938 55168
rect 42521 55165 42533 55168
rect 42567 55165 42579 55199
rect 42521 55159 42579 55165
rect 43257 55199 43315 55205
rect 43257 55165 43269 55199
rect 43303 55165 43315 55199
rect 43257 55159 43315 55165
rect 41156 55128 41184 55156
rect 42702 55128 42708 55140
rect 36279 55100 37320 55128
rect 40696 55100 42708 55128
rect 37292 55072 37320 55100
rect 42702 55088 42708 55100
rect 42760 55088 42766 55140
rect 24762 55060 24768 55072
rect 24723 55032 24768 55060
rect 24762 55020 24768 55032
rect 24820 55020 24826 55072
rect 27614 55060 27620 55072
rect 27575 55032 27620 55060
rect 27614 55020 27620 55032
rect 27672 55020 27678 55072
rect 28442 55020 28448 55072
rect 28500 55060 28506 55072
rect 28537 55063 28595 55069
rect 28537 55060 28549 55063
rect 28500 55032 28549 55060
rect 28500 55020 28506 55032
rect 28537 55029 28549 55032
rect 28583 55029 28595 55063
rect 31846 55060 31852 55072
rect 31807 55032 31852 55060
rect 28537 55023 28595 55029
rect 31846 55020 31852 55032
rect 31904 55020 31910 55072
rect 32217 55063 32275 55069
rect 32217 55029 32229 55063
rect 32263 55060 32275 55063
rect 32398 55060 32404 55072
rect 32263 55032 32404 55060
rect 32263 55029 32275 55032
rect 32217 55023 32275 55029
rect 32398 55020 32404 55032
rect 32456 55020 32462 55072
rect 37274 55020 37280 55072
rect 37332 55020 37338 55072
rect 40310 55020 40316 55072
rect 40368 55060 40374 55072
rect 40773 55063 40831 55069
rect 40773 55060 40785 55063
rect 40368 55032 40785 55060
rect 40368 55020 40374 55032
rect 40773 55029 40785 55032
rect 40819 55029 40831 55063
rect 40773 55023 40831 55029
rect 41141 55063 41199 55069
rect 41141 55029 41153 55063
rect 41187 55060 41199 55063
rect 41230 55060 41236 55072
rect 41187 55032 41236 55060
rect 41187 55029 41199 55032
rect 41141 55023 41199 55029
rect 41230 55020 41236 55032
rect 41288 55020 41294 55072
rect 41598 55060 41604 55072
rect 41559 55032 41604 55060
rect 41598 55020 41604 55032
rect 41656 55020 41662 55072
rect 41874 55060 41880 55072
rect 41835 55032 41880 55060
rect 41874 55020 41880 55032
rect 41932 55020 41938 55072
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 25777 54859 25835 54865
rect 25777 54825 25789 54859
rect 25823 54856 25835 54859
rect 26237 54859 26295 54865
rect 26237 54856 26249 54859
rect 25823 54828 26249 54856
rect 25823 54825 25835 54828
rect 25777 54819 25835 54825
rect 26237 54825 26249 54828
rect 26283 54856 26295 54859
rect 26602 54856 26608 54868
rect 26283 54828 26608 54856
rect 26283 54825 26295 54828
rect 26237 54819 26295 54825
rect 26602 54816 26608 54828
rect 26660 54816 26666 54868
rect 26694 54816 26700 54868
rect 26752 54856 26758 54868
rect 26789 54859 26847 54865
rect 26789 54856 26801 54859
rect 26752 54828 26801 54856
rect 26752 54816 26758 54828
rect 26789 54825 26801 54828
rect 26835 54825 26847 54859
rect 26789 54819 26847 54825
rect 27709 54859 27767 54865
rect 27709 54825 27721 54859
rect 27755 54856 27767 54859
rect 28074 54856 28080 54868
rect 27755 54828 28080 54856
rect 27755 54825 27767 54828
rect 27709 54819 27767 54825
rect 28074 54816 28080 54828
rect 28132 54816 28138 54868
rect 28718 54816 28724 54868
rect 28776 54856 28782 54868
rect 29089 54859 29147 54865
rect 29089 54856 29101 54859
rect 28776 54828 29101 54856
rect 28776 54816 28782 54828
rect 29089 54825 29101 54828
rect 29135 54825 29147 54859
rect 29089 54819 29147 54825
rect 29546 54816 29552 54868
rect 29604 54856 29610 54868
rect 30101 54859 30159 54865
rect 30101 54856 30113 54859
rect 29604 54828 30113 54856
rect 29604 54816 29610 54828
rect 30101 54825 30113 54828
rect 30147 54825 30159 54859
rect 30101 54819 30159 54825
rect 30834 54816 30840 54868
rect 30892 54856 30898 54868
rect 31021 54859 31079 54865
rect 31021 54856 31033 54859
rect 30892 54828 31033 54856
rect 30892 54816 30898 54828
rect 31021 54825 31033 54828
rect 31067 54825 31079 54859
rect 31021 54819 31079 54825
rect 34790 54816 34796 54868
rect 34848 54856 34854 54868
rect 35161 54859 35219 54865
rect 35161 54856 35173 54859
rect 34848 54828 35173 54856
rect 34848 54816 34854 54828
rect 35161 54825 35173 54828
rect 35207 54825 35219 54859
rect 35161 54819 35219 54825
rect 35342 54816 35348 54868
rect 35400 54856 35406 54868
rect 35805 54859 35863 54865
rect 35805 54856 35817 54859
rect 35400 54828 35817 54856
rect 35400 54816 35406 54828
rect 35805 54825 35817 54828
rect 35851 54825 35863 54859
rect 35805 54819 35863 54825
rect 36354 54816 36360 54868
rect 36412 54856 36418 54868
rect 36449 54859 36507 54865
rect 36449 54856 36461 54859
rect 36412 54828 36461 54856
rect 36412 54816 36418 54828
rect 36449 54825 36461 54828
rect 36495 54825 36507 54859
rect 36449 54819 36507 54825
rect 37185 54859 37243 54865
rect 37185 54825 37197 54859
rect 37231 54856 37243 54859
rect 37274 54856 37280 54868
rect 37231 54828 37280 54856
rect 37231 54825 37243 54828
rect 37185 54819 37243 54825
rect 37274 54816 37280 54828
rect 37332 54816 37338 54868
rect 37734 54816 37740 54868
rect 37792 54856 37798 54868
rect 37829 54859 37887 54865
rect 37829 54856 37841 54859
rect 37792 54828 37841 54856
rect 37792 54816 37798 54828
rect 37829 54825 37841 54828
rect 37875 54825 37887 54859
rect 38470 54856 38476 54868
rect 38431 54828 38476 54856
rect 37829 54819 37887 54825
rect 38470 54816 38476 54828
rect 38528 54816 38534 54868
rect 39577 54859 39635 54865
rect 39577 54825 39589 54859
rect 39623 54856 39635 54859
rect 39942 54856 39948 54868
rect 39623 54828 39948 54856
rect 39623 54825 39635 54828
rect 39577 54819 39635 54825
rect 39942 54816 39948 54828
rect 40000 54816 40006 54868
rect 41690 54856 41696 54868
rect 41651 54828 41696 54856
rect 41690 54816 41696 54828
rect 41748 54816 41754 54868
rect 44913 54859 44971 54865
rect 44913 54825 44925 54859
rect 44959 54856 44971 54859
rect 45002 54856 45008 54868
rect 44959 54828 45008 54856
rect 44959 54825 44971 54828
rect 44913 54819 44971 54825
rect 45002 54816 45008 54828
rect 45060 54816 45066 54868
rect 24397 54791 24455 54797
rect 24397 54757 24409 54791
rect 24443 54788 24455 54791
rect 24762 54788 24768 54800
rect 24443 54760 24768 54788
rect 24443 54757 24455 54760
rect 24397 54751 24455 54757
rect 24762 54748 24768 54760
rect 24820 54788 24826 54800
rect 25225 54791 25283 54797
rect 25225 54788 25237 54791
rect 24820 54760 25237 54788
rect 24820 54748 24826 54760
rect 25225 54757 25237 54760
rect 25271 54788 25283 54791
rect 26970 54788 26976 54800
rect 25271 54760 26976 54788
rect 25271 54757 25283 54760
rect 25225 54751 25283 54757
rect 26970 54748 26976 54760
rect 27028 54748 27034 54800
rect 28534 54748 28540 54800
rect 28592 54788 28598 54800
rect 28629 54791 28687 54797
rect 28629 54788 28641 54791
rect 28592 54760 28641 54788
rect 28592 54748 28598 54760
rect 28629 54757 28641 54760
rect 28675 54757 28687 54791
rect 30374 54788 30380 54800
rect 28629 54751 28687 54757
rect 29288 54760 30380 54788
rect 29288 54671 29316 54760
rect 30374 54748 30380 54760
rect 30432 54748 30438 54800
rect 39482 54788 39488 54800
rect 39316 54760 39488 54788
rect 33870 54680 33876 54732
rect 33928 54720 33934 54732
rect 35710 54720 35716 54732
rect 33928 54692 35716 54720
rect 33928 54680 33934 54692
rect 29265 54665 29323 54671
rect 28353 54655 28411 54661
rect 28353 54621 28365 54655
rect 28399 54652 28411 54655
rect 29265 54652 29277 54665
rect 28399 54631 29277 54652
rect 29311 54631 29323 54665
rect 28399 54625 29323 54631
rect 29357 54655 29415 54661
rect 28399 54624 29316 54625
rect 28399 54621 28411 54624
rect 28353 54615 28411 54621
rect 29357 54621 29369 54655
rect 29403 54621 29415 54655
rect 29534 54655 29592 54661
rect 29534 54652 29546 54655
rect 29357 54615 29415 54621
rect 29472 54624 29546 54652
rect 28629 54587 28687 54593
rect 28629 54553 28641 54587
rect 28675 54584 28687 54587
rect 29178 54584 29184 54596
rect 28675 54556 29184 54584
rect 28675 54553 28687 54556
rect 28629 54547 28687 54553
rect 29178 54544 29184 54556
rect 29236 54544 29242 54596
rect 28445 54519 28503 54525
rect 28445 54485 28457 54519
rect 28491 54516 28503 54519
rect 28994 54516 29000 54528
rect 28491 54488 29000 54516
rect 28491 54485 28503 54488
rect 28445 54479 28503 54485
rect 28994 54476 29000 54488
rect 29052 54516 29058 54528
rect 29380 54516 29408 54615
rect 29472 54528 29500 54624
rect 29534 54621 29546 54624
rect 29580 54621 29592 54655
rect 29534 54615 29592 54621
rect 29638 54612 29644 54664
rect 29696 54652 29702 54664
rect 29696 54624 29741 54652
rect 29696 54612 29702 54624
rect 30374 54612 30380 54664
rect 30432 54652 30438 54664
rect 30745 54655 30803 54661
rect 30745 54652 30757 54655
rect 30432 54624 30757 54652
rect 30432 54612 30438 54624
rect 30745 54621 30757 54624
rect 30791 54652 30803 54655
rect 31941 54655 31999 54661
rect 31941 54652 31953 54655
rect 30791 54624 31953 54652
rect 30791 54621 30803 54624
rect 30745 54615 30803 54621
rect 31941 54621 31953 54624
rect 31987 54621 31999 54655
rect 31941 54615 31999 54621
rect 32125 54655 32183 54661
rect 32125 54621 32137 54655
rect 32171 54621 32183 54655
rect 32398 54652 32404 54664
rect 32359 54624 32404 54652
rect 32125 54615 32183 54621
rect 30558 54544 30564 54596
rect 30616 54584 30622 54596
rect 30837 54587 30895 54593
rect 30837 54584 30849 54587
rect 30616 54556 30849 54584
rect 30616 54544 30622 54556
rect 30837 54553 30849 54556
rect 30883 54553 30895 54587
rect 30837 54547 30895 54553
rect 31021 54587 31079 54593
rect 31021 54553 31033 54587
rect 31067 54584 31079 54587
rect 31110 54584 31116 54596
rect 31067 54556 31116 54584
rect 31067 54553 31079 54556
rect 31021 54547 31079 54553
rect 31110 54544 31116 54556
rect 31168 54544 31174 54596
rect 32140 54584 32168 54615
rect 32398 54612 32404 54624
rect 32456 54612 32462 54664
rect 33045 54655 33103 54661
rect 33045 54621 33057 54655
rect 33091 54652 33103 54655
rect 33134 54652 33140 54664
rect 33091 54624 33140 54652
rect 33091 54621 33103 54624
rect 33045 54615 33103 54621
rect 33134 54612 33140 54624
rect 33192 54612 33198 54664
rect 33318 54652 33324 54664
rect 33279 54624 33324 54652
rect 33318 54612 33324 54624
rect 33376 54612 33382 54664
rect 34422 54652 34428 54664
rect 34383 54624 34428 54652
rect 34422 54612 34428 54624
rect 34480 54612 34486 54664
rect 34532 54661 34560 54692
rect 35710 54680 35716 54692
rect 35768 54680 35774 54732
rect 39316 54729 39344 54760
rect 39482 54748 39488 54760
rect 39540 54788 39546 54800
rect 43533 54791 43591 54797
rect 43533 54788 43545 54791
rect 39540 54760 43545 54788
rect 39540 54748 39546 54760
rect 43533 54757 43545 54760
rect 43579 54757 43591 54791
rect 43533 54751 43591 54757
rect 39301 54723 39359 54729
rect 39301 54689 39313 54723
rect 39347 54689 39359 54723
rect 39301 54683 39359 54689
rect 39850 54680 39856 54732
rect 39908 54720 39914 54732
rect 40773 54723 40831 54729
rect 40773 54720 40785 54723
rect 39908 54692 40785 54720
rect 39908 54680 39914 54692
rect 40773 54689 40785 54692
rect 40819 54720 40831 54723
rect 40862 54720 40868 54732
rect 40819 54692 40868 54720
rect 40819 54689 40831 54692
rect 40773 54683 40831 54689
rect 40862 54680 40868 54692
rect 40920 54680 40926 54732
rect 41874 54720 41880 54732
rect 40972 54692 41880 54720
rect 34517 54655 34575 54661
rect 34517 54621 34529 54655
rect 34563 54621 34575 54655
rect 34517 54615 34575 54621
rect 34606 54612 34612 54664
rect 34664 54652 34670 54664
rect 39206 54652 39212 54664
rect 34664 54624 34709 54652
rect 39167 54624 39212 54652
rect 34664 54612 34670 54624
rect 39206 54612 39212 54624
rect 39264 54612 39270 54664
rect 40972 54661 41000 54692
rect 41874 54680 41880 54692
rect 41932 54680 41938 54732
rect 43993 54723 44051 54729
rect 43993 54689 44005 54723
rect 44039 54720 44051 54723
rect 44545 54723 44603 54729
rect 44545 54720 44557 54723
rect 44039 54692 44557 54720
rect 44039 54689 44051 54692
rect 43993 54683 44051 54689
rect 44545 54689 44557 54692
rect 44591 54689 44603 54723
rect 44545 54683 44603 54689
rect 44910 54680 44916 54732
rect 44968 54720 44974 54732
rect 45005 54723 45063 54729
rect 45005 54720 45017 54723
rect 44968 54692 45017 54720
rect 44968 54680 44974 54692
rect 45005 54689 45017 54692
rect 45051 54689 45063 54723
rect 45005 54683 45063 54689
rect 40957 54655 41015 54661
rect 40957 54621 40969 54655
rect 41003 54621 41015 54655
rect 41230 54652 41236 54664
rect 41191 54624 41236 54652
rect 40957 54615 41015 54621
rect 41230 54612 41236 54624
rect 41288 54612 41294 54664
rect 42613 54655 42671 54661
rect 42613 54621 42625 54655
rect 42659 54621 42671 54655
rect 42613 54615 42671 54621
rect 32582 54584 32588 54596
rect 32140 54556 32588 54584
rect 32582 54544 32588 54556
rect 32640 54544 32646 54596
rect 38746 54544 38752 54596
rect 38804 54584 38810 54596
rect 40221 54587 40279 54593
rect 40221 54584 40233 54587
rect 38804 54556 40233 54584
rect 38804 54544 38810 54556
rect 40221 54553 40233 54556
rect 40267 54553 40279 54587
rect 40221 54547 40279 54553
rect 41141 54587 41199 54593
rect 41141 54553 41153 54587
rect 41187 54584 41199 54587
rect 41966 54584 41972 54596
rect 41187 54556 41972 54584
rect 41187 54553 41199 54556
rect 41141 54547 41199 54553
rect 41966 54544 41972 54556
rect 42024 54544 42030 54596
rect 42628 54584 42656 54615
rect 42702 54612 42708 54664
rect 42760 54652 42766 54664
rect 42760 54624 42805 54652
rect 42760 54612 42766 54624
rect 43530 54612 43536 54664
rect 43588 54652 43594 54664
rect 43901 54655 43959 54661
rect 43901 54652 43913 54655
rect 43588 54624 43913 54652
rect 43588 54612 43594 54624
rect 43901 54621 43913 54624
rect 43947 54621 43959 54655
rect 44726 54652 44732 54664
rect 44687 54624 44732 54652
rect 43901 54615 43959 54621
rect 44726 54612 44732 54624
rect 44784 54612 44790 54664
rect 44744 54584 44772 54612
rect 42628 54556 44772 54584
rect 29052 54488 29408 54516
rect 29052 54476 29058 54488
rect 29454 54476 29460 54528
rect 29512 54476 29518 54528
rect 32309 54519 32367 54525
rect 32309 54485 32321 54519
rect 32355 54516 32367 54519
rect 32858 54516 32864 54528
rect 32355 54488 32864 54516
rect 32355 54485 32367 54488
rect 32309 54479 32367 54485
rect 32858 54476 32864 54488
rect 32916 54476 32922 54528
rect 33229 54519 33287 54525
rect 33229 54485 33241 54519
rect 33275 54516 33287 54519
rect 33502 54516 33508 54528
rect 33275 54488 33508 54516
rect 33275 54485 33287 54488
rect 33229 54479 33287 54485
rect 33502 54476 33508 54488
rect 33560 54516 33566 54528
rect 34241 54519 34299 54525
rect 34241 54516 34253 54519
rect 33560 54488 34253 54516
rect 33560 54476 33566 54488
rect 34241 54485 34253 54488
rect 34287 54485 34299 54519
rect 42426 54516 42432 54528
rect 42387 54488 42432 54516
rect 34241 54479 34299 54485
rect 42426 54476 42432 54488
rect 42484 54476 42490 54528
rect 42794 54476 42800 54528
rect 42852 54516 42858 54528
rect 43073 54519 43131 54525
rect 43073 54516 43085 54519
rect 42852 54488 43085 54516
rect 42852 54476 42858 54488
rect 43073 54485 43085 54488
rect 43119 54516 43131 54519
rect 44174 54516 44180 54528
rect 43119 54488 44180 54516
rect 43119 54485 43131 54488
rect 43073 54479 43131 54485
rect 44174 54476 44180 54488
rect 44232 54476 44238 54528
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 27062 54272 27068 54324
rect 27120 54312 27126 54324
rect 27249 54315 27307 54321
rect 27249 54312 27261 54315
rect 27120 54284 27261 54312
rect 27120 54272 27126 54284
rect 27249 54281 27261 54284
rect 27295 54281 27307 54315
rect 27890 54312 27896 54324
rect 27851 54284 27896 54312
rect 27249 54275 27307 54281
rect 27890 54272 27896 54284
rect 27948 54272 27954 54324
rect 28902 54312 28908 54324
rect 28863 54284 28908 54312
rect 28902 54272 28908 54284
rect 28960 54272 28966 54324
rect 29178 54272 29184 54324
rect 29236 54312 29242 54324
rect 29365 54315 29423 54321
rect 29365 54312 29377 54315
rect 29236 54284 29377 54312
rect 29236 54272 29242 54284
rect 29365 54281 29377 54284
rect 29411 54312 29423 54315
rect 29638 54312 29644 54324
rect 29411 54284 29644 54312
rect 29411 54281 29423 54284
rect 29365 54275 29423 54281
rect 29638 54272 29644 54284
rect 29696 54272 29702 54324
rect 32769 54315 32827 54321
rect 32769 54281 32781 54315
rect 32815 54312 32827 54315
rect 33226 54312 33232 54324
rect 32815 54284 33232 54312
rect 32815 54281 32827 54284
rect 32769 54275 32827 54281
rect 33226 54272 33232 54284
rect 33284 54272 33290 54324
rect 33318 54272 33324 54324
rect 33376 54312 33382 54324
rect 33597 54315 33655 54321
rect 33597 54312 33609 54315
rect 33376 54284 33609 54312
rect 33376 54272 33382 54284
rect 33597 54281 33609 54284
rect 33643 54281 33655 54315
rect 33597 54275 33655 54281
rect 34241 54315 34299 54321
rect 34241 54281 34253 54315
rect 34287 54312 34299 54315
rect 34606 54312 34612 54324
rect 34287 54284 34612 54312
rect 34287 54281 34299 54284
rect 34241 54275 34299 54281
rect 34606 54272 34612 54284
rect 34664 54272 34670 54324
rect 34974 54272 34980 54324
rect 35032 54312 35038 54324
rect 35434 54312 35440 54324
rect 35032 54284 35440 54312
rect 35032 54272 35038 54284
rect 35434 54272 35440 54284
rect 35492 54272 35498 54324
rect 36446 54272 36452 54324
rect 36504 54312 36510 54324
rect 36633 54315 36691 54321
rect 36633 54312 36645 54315
rect 36504 54284 36645 54312
rect 36504 54272 36510 54284
rect 36633 54281 36645 54284
rect 36679 54281 36691 54315
rect 36633 54275 36691 54281
rect 37182 54272 37188 54324
rect 37240 54312 37246 54324
rect 37277 54315 37335 54321
rect 37277 54312 37289 54315
rect 37240 54284 37289 54312
rect 37240 54272 37246 54284
rect 37277 54281 37289 54284
rect 37323 54281 37335 54315
rect 39022 54312 39028 54324
rect 38983 54284 39028 54312
rect 37277 54275 37335 54281
rect 39022 54272 39028 54284
rect 39080 54272 39086 54324
rect 40310 54312 40316 54324
rect 40271 54284 40316 54312
rect 40310 54272 40316 54284
rect 40368 54272 40374 54324
rect 41414 54272 41420 54324
rect 41472 54312 41478 54324
rect 41509 54315 41567 54321
rect 41509 54312 41521 54315
rect 41472 54284 41521 54312
rect 41472 54272 41478 54284
rect 41509 54281 41521 54284
rect 41555 54281 41567 54315
rect 41966 54312 41972 54324
rect 41927 54284 41972 54312
rect 41509 54275 41567 54281
rect 41966 54272 41972 54284
rect 42024 54272 42030 54324
rect 29730 54204 29736 54256
rect 29788 54244 29794 54256
rect 32674 54244 32680 54256
rect 29788 54216 32680 54244
rect 29788 54204 29794 54216
rect 28534 54176 28540 54188
rect 28495 54148 28540 54176
rect 28534 54136 28540 54148
rect 28592 54136 28598 54188
rect 30392 54185 30420 54216
rect 32674 54204 32680 54216
rect 32732 54204 32738 54256
rect 39669 54247 39727 54253
rect 34440 54216 36032 54244
rect 34440 54188 34468 54216
rect 29549 54179 29607 54185
rect 29549 54145 29561 54179
rect 29595 54176 29607 54179
rect 30377 54179 30435 54185
rect 29595 54148 30236 54176
rect 29595 54145 29607 54148
rect 29549 54139 29607 54145
rect 28442 54108 28448 54120
rect 28403 54080 28448 54108
rect 28442 54068 28448 54080
rect 28500 54068 28506 54120
rect 29730 54108 29736 54120
rect 29691 54080 29736 54108
rect 29730 54068 29736 54080
rect 29788 54068 29794 54120
rect 30208 54052 30236 54148
rect 30377 54145 30389 54179
rect 30423 54145 30435 54179
rect 32398 54176 32404 54188
rect 32359 54148 32404 54176
rect 30377 54139 30435 54145
rect 32398 54136 32404 54148
rect 32456 54136 32462 54188
rect 33781 54179 33839 54185
rect 33781 54145 33793 54179
rect 33827 54176 33839 54179
rect 34422 54176 34428 54188
rect 33827 54148 34428 54176
rect 33827 54145 33839 54148
rect 33781 54139 33839 54145
rect 34422 54136 34428 54148
rect 34480 54136 34486 54188
rect 34974 54136 34980 54188
rect 35032 54185 35038 54188
rect 35032 54179 35049 54185
rect 35037 54145 35049 54179
rect 35710 54176 35716 54188
rect 35671 54148 35716 54176
rect 35032 54139 35049 54145
rect 35032 54136 35038 54139
rect 35710 54136 35716 54148
rect 35768 54136 35774 54188
rect 36004 54185 36032 54216
rect 39669 54213 39681 54247
rect 39715 54244 39727 54247
rect 40218 54244 40224 54256
rect 39715 54216 40224 54244
rect 39715 54213 39727 54216
rect 39669 54207 39727 54213
rect 35989 54179 36047 54185
rect 35989 54145 36001 54179
rect 36035 54145 36047 54179
rect 35989 54139 36047 54145
rect 38194 54136 38200 54188
rect 38252 54176 38258 54188
rect 38289 54179 38347 54185
rect 38289 54176 38301 54179
rect 38252 54148 38301 54176
rect 38252 54136 38258 54148
rect 38289 54145 38301 54148
rect 38335 54145 38347 54179
rect 38289 54139 38347 54145
rect 39117 54179 39175 54185
rect 39117 54145 39129 54179
rect 39163 54176 39175 54179
rect 39684 54176 39712 54207
rect 40218 54204 40224 54216
rect 40276 54204 40282 54256
rect 42058 54204 42064 54256
rect 42116 54244 42122 54256
rect 42337 54247 42395 54253
rect 42337 54244 42349 54247
rect 42116 54216 42349 54244
rect 42116 54204 42122 54216
rect 42337 54213 42349 54216
rect 42383 54244 42395 54247
rect 43257 54247 43315 54253
rect 43257 54244 43269 54247
rect 42383 54216 43269 54244
rect 42383 54213 42395 54216
rect 42337 54207 42395 54213
rect 43257 54213 43269 54216
rect 43303 54213 43315 54247
rect 44726 54244 44732 54256
rect 43257 54207 43315 54213
rect 43456 54216 44732 54244
rect 39163 54148 39712 54176
rect 39163 54145 39175 54148
rect 39117 54139 39175 54145
rect 40034 54136 40040 54188
rect 40092 54176 40098 54188
rect 40129 54179 40187 54185
rect 40129 54176 40141 54179
rect 40092 54148 40141 54176
rect 40092 54136 40098 54148
rect 40129 54145 40141 54148
rect 40175 54145 40187 54179
rect 40129 54139 40187 54145
rect 41141 54179 41199 54185
rect 41141 54145 41153 54179
rect 41187 54176 41199 54179
rect 41598 54176 41604 54188
rect 41187 54148 41604 54176
rect 41187 54145 41199 54148
rect 41141 54139 41199 54145
rect 41598 54136 41604 54148
rect 41656 54136 41662 54188
rect 42153 54179 42211 54185
rect 42153 54145 42165 54179
rect 42199 54145 42211 54179
rect 42426 54176 42432 54188
rect 42387 54148 42432 54176
rect 42153 54139 42211 54145
rect 30469 54111 30527 54117
rect 30469 54077 30481 54111
rect 30515 54077 30527 54111
rect 30469 54071 30527 54077
rect 26605 54043 26663 54049
rect 26605 54009 26617 54043
rect 26651 54040 26663 54043
rect 26970 54040 26976 54052
rect 26651 54012 26976 54040
rect 26651 54009 26663 54012
rect 26605 54003 26663 54009
rect 26970 54000 26976 54012
rect 27028 54040 27034 54052
rect 28626 54040 28632 54052
rect 27028 54012 28632 54040
rect 27028 54000 27034 54012
rect 28626 54000 28632 54012
rect 28684 54000 28690 54052
rect 30190 54000 30196 54052
rect 30248 54040 30254 54052
rect 30484 54040 30512 54071
rect 30558 54068 30564 54120
rect 30616 54108 30622 54120
rect 30745 54111 30803 54117
rect 30745 54108 30757 54111
rect 30616 54080 30757 54108
rect 30616 54068 30622 54080
rect 30745 54077 30757 54080
rect 30791 54077 30803 54111
rect 32306 54108 32312 54120
rect 32267 54080 32312 54108
rect 30745 54071 30803 54077
rect 32306 54068 32312 54080
rect 32364 54068 32370 54120
rect 33870 54108 33876 54120
rect 33831 54080 33876 54108
rect 33870 54068 33876 54080
rect 33928 54068 33934 54120
rect 35161 54111 35219 54117
rect 35161 54077 35173 54111
rect 35207 54077 35219 54111
rect 41230 54108 41236 54120
rect 41191 54080 41236 54108
rect 35161 54071 35219 54077
rect 34701 54043 34759 54049
rect 34701 54040 34713 54043
rect 30248 54012 34713 54040
rect 30248 54000 30254 54012
rect 34701 54009 34713 54012
rect 34747 54009 34759 54043
rect 35176 54040 35204 54071
rect 41230 54068 41236 54080
rect 41288 54068 41294 54120
rect 42168 54108 42196 54139
rect 42426 54136 42432 54148
rect 42484 54136 42490 54188
rect 43456 54185 43484 54216
rect 44726 54204 44732 54216
rect 44784 54204 44790 54256
rect 43441 54179 43499 54185
rect 43441 54145 43453 54179
rect 43487 54145 43499 54179
rect 43441 54139 43499 54145
rect 43533 54179 43591 54185
rect 43533 54145 43545 54179
rect 43579 54145 43591 54179
rect 43533 54139 43591 54145
rect 43625 54179 43683 54185
rect 43625 54145 43637 54179
rect 43671 54176 43683 54179
rect 44174 54176 44180 54188
rect 43671 54148 44180 54176
rect 43671 54145 43683 54148
rect 43625 54139 43683 54145
rect 42242 54108 42248 54120
rect 42155 54080 42248 54108
rect 42242 54068 42248 54080
rect 42300 54108 42306 54120
rect 42610 54108 42616 54120
rect 42300 54080 42616 54108
rect 42300 54068 42306 54080
rect 42610 54068 42616 54080
rect 42668 54068 42674 54120
rect 42702 54068 42708 54120
rect 42760 54108 42766 54120
rect 43548 54108 43576 54139
rect 44174 54136 44180 54148
rect 44232 54176 44238 54188
rect 45002 54176 45008 54188
rect 44232 54148 45008 54176
rect 44232 54136 44238 54148
rect 45002 54136 45008 54148
rect 45060 54136 45066 54188
rect 44910 54108 44916 54120
rect 42760 54080 44916 54108
rect 42760 54068 42766 54080
rect 44910 54068 44916 54080
rect 44968 54068 44974 54120
rect 36173 54043 36231 54049
rect 36173 54040 36185 54043
rect 35176 54012 36185 54040
rect 34701 54003 34759 54009
rect 36173 54009 36185 54012
rect 36219 54009 36231 54043
rect 36173 54003 36231 54009
rect 31110 53932 31116 53984
rect 31168 53972 31174 53984
rect 31389 53975 31447 53981
rect 31389 53972 31401 53975
rect 31168 53944 31401 53972
rect 31168 53932 31174 53944
rect 31389 53941 31401 53944
rect 31435 53972 31447 53975
rect 33686 53972 33692 53984
rect 31435 53944 33692 53972
rect 31435 53941 31447 53944
rect 31389 53935 31447 53941
rect 33686 53932 33692 53944
rect 33744 53932 33750 53984
rect 34606 53932 34612 53984
rect 34664 53972 34670 53984
rect 35805 53975 35863 53981
rect 35805 53972 35817 53975
rect 34664 53944 35817 53972
rect 34664 53932 34670 53944
rect 35805 53941 35817 53944
rect 35851 53941 35863 53975
rect 35805 53935 35863 53941
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 28994 53728 29000 53780
rect 29052 53768 29058 53780
rect 29825 53771 29883 53777
rect 29825 53768 29837 53771
rect 29052 53740 29837 53768
rect 29052 53728 29058 53740
rect 29825 53737 29837 53740
rect 29871 53737 29883 53771
rect 32398 53768 32404 53780
rect 32359 53740 32404 53768
rect 29825 53731 29883 53737
rect 32398 53728 32404 53740
rect 32456 53728 32462 53780
rect 32582 53768 32588 53780
rect 32543 53740 32588 53768
rect 32582 53728 32588 53740
rect 32640 53768 32646 53780
rect 33321 53771 33379 53777
rect 33321 53768 33333 53771
rect 32640 53740 33333 53768
rect 32640 53728 32646 53740
rect 33321 53737 33333 53740
rect 33367 53737 33379 53771
rect 33502 53768 33508 53780
rect 33463 53740 33508 53768
rect 33321 53731 33379 53737
rect 33502 53728 33508 53740
rect 33560 53728 33566 53780
rect 34882 53768 34888 53780
rect 34795 53740 34888 53768
rect 34882 53728 34888 53740
rect 34940 53768 34946 53780
rect 35437 53771 35495 53777
rect 35437 53768 35449 53771
rect 34940 53740 35449 53768
rect 34940 53728 34946 53740
rect 35437 53737 35449 53740
rect 35483 53768 35495 53771
rect 35526 53768 35532 53780
rect 35483 53740 35532 53768
rect 35483 53737 35495 53740
rect 35437 53731 35495 53737
rect 35526 53728 35532 53740
rect 35584 53728 35590 53780
rect 35894 53768 35900 53780
rect 35855 53740 35900 53768
rect 35894 53728 35900 53740
rect 35952 53728 35958 53780
rect 40034 53728 40040 53780
rect 40092 53768 40098 53780
rect 40221 53771 40279 53777
rect 40221 53768 40233 53771
rect 40092 53740 40233 53768
rect 40092 53728 40098 53740
rect 40221 53737 40233 53740
rect 40267 53737 40279 53771
rect 41874 53768 41880 53780
rect 41835 53740 41880 53768
rect 40221 53731 40279 53737
rect 41874 53728 41880 53740
rect 41932 53728 41938 53780
rect 42058 53768 42064 53780
rect 42019 53740 42064 53768
rect 42058 53728 42064 53740
rect 42116 53728 42122 53780
rect 27525 53703 27583 53709
rect 27525 53669 27537 53703
rect 27571 53700 27583 53703
rect 29181 53703 29239 53709
rect 29181 53700 29193 53703
rect 27571 53672 29193 53700
rect 27571 53669 27583 53672
rect 27525 53663 27583 53669
rect 29181 53669 29193 53672
rect 29227 53700 29239 53703
rect 31110 53700 31116 53712
rect 29227 53672 31116 53700
rect 29227 53669 29239 53672
rect 29181 53663 29239 53669
rect 31110 53660 31116 53672
rect 31168 53660 31174 53712
rect 33686 53660 33692 53712
rect 33744 53700 33750 53712
rect 34333 53703 34391 53709
rect 34333 53700 34345 53703
rect 33744 53672 34345 53700
rect 33744 53660 33750 53672
rect 34333 53669 34345 53672
rect 34379 53700 34391 53703
rect 36446 53700 36452 53712
rect 34379 53672 36452 53700
rect 34379 53669 34391 53672
rect 34333 53663 34391 53669
rect 36446 53660 36452 53672
rect 36504 53660 36510 53712
rect 33134 53592 33140 53644
rect 33192 53632 33198 53644
rect 33192 53604 33732 53632
rect 33192 53592 33198 53604
rect 29730 53524 29736 53576
rect 29788 53564 29794 53576
rect 30009 53567 30067 53573
rect 30009 53564 30021 53567
rect 29788 53536 30021 53564
rect 29788 53524 29794 53536
rect 30009 53533 30021 53536
rect 30055 53533 30067 53567
rect 30190 53564 30196 53576
rect 30151 53536 30196 53564
rect 30009 53527 30067 53533
rect 30190 53524 30196 53536
rect 30248 53524 30254 53576
rect 32858 53564 32864 53576
rect 32819 53536 32864 53564
rect 32858 53524 32864 53536
rect 32916 53524 32922 53576
rect 33318 53524 33324 53576
rect 33376 53524 33382 53576
rect 33336 53496 33364 53524
rect 33704 53505 33732 53604
rect 40218 53592 40224 53644
rect 40276 53632 40282 53644
rect 40770 53632 40776 53644
rect 40276 53604 40776 53632
rect 40276 53592 40282 53604
rect 40770 53592 40776 53604
rect 40828 53632 40834 53644
rect 41325 53635 41383 53641
rect 41325 53632 41337 53635
rect 40828 53604 41337 53632
rect 40828 53592 40834 53604
rect 41325 53601 41337 53604
rect 41371 53601 41383 53635
rect 41325 53595 41383 53601
rect 33473 53499 33531 53505
rect 33473 53496 33485 53499
rect 33336 53468 33485 53496
rect 33473 53465 33485 53468
rect 33519 53465 33531 53499
rect 33473 53459 33531 53465
rect 33689 53499 33747 53505
rect 33689 53465 33701 53499
rect 33735 53465 33747 53499
rect 42242 53496 42248 53508
rect 42203 53468 42248 53496
rect 33689 53459 33747 53465
rect 42242 53456 42248 53468
rect 42300 53456 42306 53508
rect 28626 53428 28632 53440
rect 28539 53400 28632 53428
rect 28626 53388 28632 53400
rect 28684 53428 28690 53440
rect 28994 53428 29000 53440
rect 28684 53400 29000 53428
rect 28684 53388 28690 53400
rect 28994 53388 29000 53400
rect 29052 53388 29058 53440
rect 42045 53431 42103 53437
rect 42045 53397 42057 53431
rect 42091 53428 42103 53431
rect 42426 53428 42432 53440
rect 42091 53400 42432 53428
rect 42091 53397 42103 53400
rect 42045 53391 42103 53397
rect 42426 53388 42432 53400
rect 42484 53388 42490 53440
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 33686 53224 33692 53236
rect 33647 53196 33692 53224
rect 33686 53184 33692 53196
rect 33744 53184 33750 53236
rect 34698 53184 34704 53236
rect 34756 53224 34762 53236
rect 35345 53227 35403 53233
rect 35345 53224 35357 53227
rect 34756 53196 35357 53224
rect 34756 53184 34762 53196
rect 35345 53193 35357 53196
rect 35391 53193 35403 53227
rect 40770 53224 40776 53236
rect 40731 53196 40776 53224
rect 35345 53187 35403 53193
rect 40770 53184 40776 53196
rect 40828 53184 40834 53236
rect 32585 53159 32643 53165
rect 32585 53125 32597 53159
rect 32631 53156 32643 53159
rect 33229 53159 33287 53165
rect 33229 53156 33241 53159
rect 32631 53128 33241 53156
rect 32631 53125 32643 53128
rect 32585 53119 32643 53125
rect 33229 53125 33241 53128
rect 33275 53156 33287 53159
rect 34333 53159 34391 53165
rect 34333 53156 34345 53159
rect 33275 53128 34345 53156
rect 33275 53125 33287 53128
rect 33229 53119 33287 53125
rect 34333 53125 34345 53128
rect 34379 53156 34391 53159
rect 34882 53156 34888 53168
rect 34379 53128 34888 53156
rect 34379 53125 34391 53128
rect 34333 53119 34391 53125
rect 34882 53116 34888 53128
rect 34940 53116 34946 53168
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 27522 52368 27528 52420
rect 27580 52408 27586 52420
rect 34514 52408 34520 52420
rect 27580 52380 34520 52408
rect 27580 52368 27586 52380
rect 34514 52368 34520 52380
rect 34572 52368 34578 52420
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 34241 52071 34299 52077
rect 34241 52037 34253 52071
rect 34287 52068 34299 52071
rect 34514 52068 34520 52080
rect 34287 52040 34520 52068
rect 34287 52037 34299 52040
rect 34241 52031 34299 52037
rect 34514 52028 34520 52040
rect 34572 52028 34578 52080
rect 34054 51932 34060 51944
rect 34015 51904 34060 51932
rect 34054 51892 34060 51904
rect 34112 51892 34118 51944
rect 35802 51932 35808 51944
rect 35763 51904 35808 51932
rect 35802 51892 35808 51904
rect 35860 51892 35866 51944
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 34054 51552 34060 51604
rect 34112 51592 34118 51604
rect 34241 51595 34299 51601
rect 34241 51592 34253 51595
rect 34112 51564 34253 51592
rect 34112 51552 34118 51564
rect 34241 51561 34253 51564
rect 34287 51561 34299 51595
rect 34241 51555 34299 51561
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 29546 8440 29552 8492
rect 29604 8480 29610 8492
rect 30009 8483 30067 8489
rect 30009 8480 30021 8483
rect 29604 8452 30021 8480
rect 29604 8440 29610 8452
rect 30009 8449 30021 8452
rect 30055 8449 30067 8483
rect 30009 8443 30067 8449
rect 30101 8347 30159 8353
rect 30101 8313 30113 8347
rect 30147 8344 30159 8347
rect 30190 8344 30196 8356
rect 30147 8316 30196 8344
rect 30147 8313 30159 8316
rect 30101 8307 30159 8313
rect 30190 8304 30196 8316
rect 30248 8304 30254 8356
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 28994 8072 29000 8084
rect 28955 8044 29000 8072
rect 28994 8032 29000 8044
rect 29052 8032 29058 8084
rect 29546 7896 29552 7948
rect 29604 7936 29610 7948
rect 29604 7908 30880 7936
rect 29604 7896 29610 7908
rect 29454 7868 29460 7880
rect 29415 7840 29460 7868
rect 29454 7828 29460 7840
rect 29512 7828 29518 7880
rect 30006 7828 30012 7880
rect 30064 7868 30070 7880
rect 30852 7877 30880 7908
rect 30101 7871 30159 7877
rect 30101 7868 30113 7871
rect 30064 7840 30113 7868
rect 30064 7828 30070 7840
rect 30101 7837 30113 7840
rect 30147 7837 30159 7871
rect 30101 7831 30159 7837
rect 30837 7871 30895 7877
rect 30837 7837 30849 7871
rect 30883 7837 30895 7871
rect 30837 7831 30895 7837
rect 30929 7735 30987 7741
rect 30929 7701 30941 7735
rect 30975 7732 30987 7735
rect 31202 7732 31208 7744
rect 30975 7704 31208 7732
rect 30975 7701 30987 7704
rect 30929 7695 30987 7701
rect 31202 7692 31208 7704
rect 31260 7692 31266 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 26970 7392 26976 7404
rect 26931 7364 26976 7392
rect 26970 7352 26976 7364
rect 27028 7352 27034 7404
rect 29086 7352 29092 7404
rect 29144 7392 29150 7404
rect 30009 7395 30067 7401
rect 30009 7392 30021 7395
rect 29144 7364 30021 7392
rect 29144 7352 29150 7364
rect 30009 7361 30021 7364
rect 30055 7361 30067 7395
rect 30009 7355 30067 7361
rect 31570 7352 31576 7404
rect 31628 7392 31634 7404
rect 32125 7395 32183 7401
rect 32125 7392 32137 7395
rect 31628 7364 32137 7392
rect 31628 7352 31634 7364
rect 32125 7361 32137 7364
rect 32171 7361 32183 7395
rect 32125 7355 32183 7361
rect 27706 7324 27712 7336
rect 27667 7296 27712 7324
rect 27706 7284 27712 7296
rect 27764 7284 27770 7336
rect 27890 7324 27896 7336
rect 27851 7296 27896 7324
rect 27890 7284 27896 7296
rect 27948 7284 27954 7336
rect 29178 7324 29184 7336
rect 29139 7296 29184 7324
rect 29178 7284 29184 7296
rect 29236 7284 29242 7336
rect 29546 7284 29552 7336
rect 29604 7324 29610 7336
rect 30193 7327 30251 7333
rect 30193 7324 30205 7327
rect 29604 7296 30205 7324
rect 29604 7284 29610 7296
rect 30193 7293 30205 7296
rect 30239 7293 30251 7327
rect 30193 7287 30251 7293
rect 26878 7188 26884 7200
rect 26839 7160 26884 7188
rect 26878 7148 26884 7160
rect 26936 7148 26942 7200
rect 31294 7188 31300 7200
rect 31255 7160 31300 7188
rect 31294 7148 31300 7160
rect 31352 7148 31358 7200
rect 32217 7191 32275 7197
rect 32217 7157 32229 7191
rect 32263 7188 32275 7191
rect 33778 7188 33784 7200
rect 32263 7160 33784 7188
rect 32263 7157 32275 7160
rect 32217 7151 32275 7157
rect 33778 7148 33784 7160
rect 33836 7148 33842 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 30558 6944 30564 6996
rect 30616 6984 30622 6996
rect 31570 6984 31576 6996
rect 30616 6956 31576 6984
rect 30616 6944 30622 6956
rect 31570 6944 31576 6956
rect 31628 6944 31634 6996
rect 28721 6851 28779 6857
rect 28721 6817 28733 6851
rect 28767 6848 28779 6851
rect 29454 6848 29460 6860
rect 28767 6820 29460 6848
rect 28767 6817 28779 6820
rect 28721 6811 28779 6817
rect 29454 6808 29460 6820
rect 29512 6808 29518 6860
rect 30282 6848 30288 6860
rect 30243 6820 30288 6848
rect 30282 6808 30288 6820
rect 30340 6808 30346 6860
rect 31202 6848 31208 6860
rect 31163 6820 31208 6848
rect 31202 6808 31208 6820
rect 31260 6808 31266 6860
rect 31478 6848 31484 6860
rect 31439 6820 31484 6848
rect 31478 6808 31484 6820
rect 31536 6808 31542 6860
rect 31570 6808 31576 6860
rect 31628 6848 31634 6860
rect 31628 6820 34284 6848
rect 31628 6808 31634 6820
rect 26881 6783 26939 6789
rect 26881 6749 26893 6783
rect 26927 6780 26939 6783
rect 26970 6780 26976 6792
rect 26927 6752 26976 6780
rect 26927 6749 26939 6752
rect 26881 6743 26939 6749
rect 26970 6740 26976 6752
rect 27028 6740 27034 6792
rect 27614 6740 27620 6792
rect 27672 6780 27678 6792
rect 34256 6789 34284 6820
rect 27709 6783 27767 6789
rect 27709 6780 27721 6783
rect 27672 6752 27721 6780
rect 27672 6740 27678 6752
rect 27709 6749 27721 6752
rect 27755 6749 27767 6783
rect 27709 6743 27767 6749
rect 31021 6783 31079 6789
rect 31021 6749 31033 6783
rect 31067 6749 31079 6783
rect 31021 6743 31079 6749
rect 34241 6783 34299 6789
rect 34241 6749 34253 6783
rect 34287 6749 34299 6783
rect 34241 6743 34299 6749
rect 28905 6715 28963 6721
rect 28905 6681 28917 6715
rect 28951 6712 28963 6715
rect 29454 6712 29460 6724
rect 28951 6684 29460 6712
rect 28951 6681 28963 6684
rect 28905 6675 28963 6681
rect 29454 6672 29460 6684
rect 29512 6672 29518 6724
rect 31036 6712 31064 6743
rect 31294 6712 31300 6724
rect 31036 6684 31300 6712
rect 31294 6672 31300 6684
rect 31352 6672 31358 6724
rect 26418 6644 26424 6656
rect 26379 6616 26424 6644
rect 26418 6604 26424 6616
rect 26476 6604 26482 6656
rect 26973 6647 27031 6653
rect 26973 6613 26985 6647
rect 27019 6644 27031 6647
rect 27798 6644 27804 6656
rect 27019 6616 27804 6644
rect 27019 6613 27031 6616
rect 26973 6607 27031 6613
rect 27798 6604 27804 6616
rect 27856 6604 27862 6656
rect 34333 6647 34391 6653
rect 34333 6613 34345 6647
rect 34379 6644 34391 6647
rect 34422 6644 34428 6656
rect 34379 6616 34428 6644
rect 34379 6613 34391 6616
rect 34333 6607 34391 6613
rect 34422 6604 34428 6616
rect 34480 6604 34486 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 29086 6440 29092 6452
rect 27448 6412 29092 6440
rect 26418 6264 26424 6316
rect 26476 6304 26482 6316
rect 26697 6307 26755 6313
rect 26697 6304 26709 6307
rect 26476 6276 26709 6304
rect 26476 6264 26482 6276
rect 26697 6273 26709 6276
rect 26743 6304 26755 6307
rect 27448 6304 27476 6412
rect 29086 6400 29092 6412
rect 29144 6400 29150 6452
rect 27798 6372 27804 6384
rect 27759 6344 27804 6372
rect 27798 6332 27804 6344
rect 27856 6332 27862 6384
rect 30558 6372 30564 6384
rect 30519 6344 30564 6372
rect 30558 6332 30564 6344
rect 30616 6332 30622 6384
rect 27614 6304 27620 6316
rect 26743 6276 27476 6304
rect 27575 6276 27620 6304
rect 26743 6273 26755 6276
rect 26697 6267 26755 6273
rect 27614 6264 27620 6276
rect 27672 6264 27678 6316
rect 29086 6264 29092 6316
rect 29144 6304 29150 6316
rect 30285 6307 30343 6313
rect 30285 6304 30297 6307
rect 29144 6276 30297 6304
rect 29144 6264 29150 6276
rect 30285 6273 30297 6276
rect 30331 6304 30343 6307
rect 31297 6307 31355 6313
rect 31297 6304 31309 6307
rect 30331 6276 31309 6304
rect 30331 6273 30343 6276
rect 30285 6267 30343 6273
rect 31297 6273 31309 6276
rect 31343 6273 31355 6307
rect 31297 6267 31355 6273
rect 26970 6236 26976 6248
rect 26883 6208 26976 6236
rect 26970 6196 26976 6208
rect 27028 6236 27034 6248
rect 27430 6236 27436 6248
rect 27028 6208 27436 6236
rect 27028 6196 27034 6208
rect 27430 6196 27436 6208
rect 27488 6196 27494 6248
rect 28074 6236 28080 6248
rect 28035 6208 28080 6236
rect 28074 6196 28080 6208
rect 28132 6196 28138 6248
rect 32582 6236 32588 6248
rect 32543 6208 32588 6236
rect 32582 6196 32588 6208
rect 32640 6196 32646 6248
rect 33042 6196 33048 6248
rect 33100 6236 33106 6248
rect 33505 6239 33563 6245
rect 33505 6236 33517 6239
rect 33100 6208 33517 6236
rect 33100 6196 33106 6208
rect 33505 6205 33517 6208
rect 33551 6205 33563 6239
rect 33505 6199 33563 6205
rect 33689 6239 33747 6245
rect 33689 6205 33701 6239
rect 33735 6205 33747 6239
rect 33689 6199 33747 6205
rect 26237 6171 26295 6177
rect 26237 6137 26249 6171
rect 26283 6168 26295 6171
rect 27706 6168 27712 6180
rect 26283 6140 27712 6168
rect 26283 6137 26295 6140
rect 26237 6131 26295 6137
rect 27706 6128 27712 6140
rect 27764 6128 27770 6180
rect 32490 6128 32496 6180
rect 32548 6168 32554 6180
rect 33704 6168 33732 6199
rect 32548 6140 33732 6168
rect 32548 6128 32554 6140
rect 25314 6100 25320 6112
rect 25275 6072 25320 6100
rect 25314 6060 25320 6072
rect 25372 6060 25378 6112
rect 34238 6060 34244 6112
rect 34296 6100 34302 6112
rect 34333 6103 34391 6109
rect 34333 6100 34345 6103
rect 34296 6072 34345 6100
rect 34296 6060 34302 6072
rect 34333 6069 34345 6072
rect 34379 6069 34391 6103
rect 34333 6063 34391 6069
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 29454 5896 29460 5908
rect 29415 5868 29460 5896
rect 29454 5856 29460 5868
rect 29512 5856 29518 5908
rect 32490 5896 32496 5908
rect 32451 5868 32496 5896
rect 32490 5856 32496 5868
rect 32548 5856 32554 5908
rect 33042 5896 33048 5908
rect 33003 5868 33048 5896
rect 33042 5856 33048 5868
rect 33100 5856 33106 5908
rect 26418 5828 26424 5840
rect 24596 5800 26424 5828
rect 24596 5701 24624 5800
rect 26418 5788 26424 5800
rect 26476 5788 26482 5840
rect 33870 5788 33876 5840
rect 33928 5828 33934 5840
rect 33928 5800 34744 5828
rect 33928 5788 33934 5800
rect 26053 5763 26111 5769
rect 26053 5729 26065 5763
rect 26099 5760 26111 5763
rect 26878 5760 26884 5772
rect 26099 5732 26884 5760
rect 26099 5729 26111 5732
rect 26053 5723 26111 5729
rect 26878 5720 26884 5732
rect 26936 5720 26942 5772
rect 27522 5760 27528 5772
rect 27483 5732 27528 5760
rect 27522 5720 27528 5732
rect 27580 5720 27586 5772
rect 30006 5760 30012 5772
rect 29967 5732 30012 5760
rect 30006 5720 30012 5732
rect 30064 5720 30070 5772
rect 30190 5760 30196 5772
rect 30151 5732 30196 5760
rect 30190 5720 30196 5732
rect 30248 5720 30254 5772
rect 30558 5760 30564 5772
rect 30519 5732 30564 5760
rect 30558 5720 30564 5732
rect 30616 5720 30622 5772
rect 30650 5720 30656 5772
rect 30708 5760 30714 5772
rect 34238 5760 34244 5772
rect 30708 5732 32996 5760
rect 34199 5732 34244 5760
rect 30708 5720 30714 5732
rect 24121 5695 24179 5701
rect 24121 5661 24133 5695
rect 24167 5692 24179 5695
rect 24581 5695 24639 5701
rect 24581 5692 24593 5695
rect 24167 5664 24593 5692
rect 24167 5661 24179 5664
rect 24121 5655 24179 5661
rect 24581 5661 24593 5664
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 25409 5695 25467 5701
rect 25409 5661 25421 5695
rect 25455 5692 25467 5695
rect 25869 5695 25927 5701
rect 25869 5692 25881 5695
rect 25455 5664 25881 5692
rect 25455 5661 25467 5664
rect 25409 5655 25467 5661
rect 25869 5661 25881 5664
rect 25915 5661 25927 5695
rect 28902 5692 28908 5704
rect 28863 5664 28908 5692
rect 25869 5655 25927 5661
rect 28902 5652 28908 5664
rect 28960 5652 28966 5704
rect 28994 5652 29000 5704
rect 29052 5692 29058 5704
rect 29546 5692 29552 5704
rect 29052 5664 29552 5692
rect 29052 5652 29058 5664
rect 29546 5652 29552 5664
rect 29604 5652 29610 5704
rect 32968 5701 32996 5732
rect 34238 5720 34244 5732
rect 34296 5720 34302 5772
rect 34422 5760 34428 5772
rect 34383 5732 34428 5760
rect 34422 5720 34428 5732
rect 34480 5720 34486 5772
rect 34716 5769 34744 5800
rect 34701 5763 34759 5769
rect 34701 5729 34713 5763
rect 34747 5729 34759 5763
rect 34701 5723 34759 5729
rect 32953 5695 33011 5701
rect 32953 5661 32965 5695
rect 32999 5661 33011 5695
rect 32953 5655 33011 5661
rect 24673 5559 24731 5565
rect 24673 5525 24685 5559
rect 24719 5556 24731 5559
rect 25498 5556 25504 5568
rect 24719 5528 25504 5556
rect 24719 5525 24731 5528
rect 24673 5519 24731 5525
rect 25498 5516 25504 5528
rect 25556 5516 25562 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 27709 5355 27767 5361
rect 27709 5321 27721 5355
rect 27755 5352 27767 5355
rect 27890 5352 27896 5364
rect 27755 5324 27896 5352
rect 27755 5321 27767 5324
rect 27709 5315 27767 5321
rect 27890 5312 27896 5324
rect 27948 5312 27954 5364
rect 25498 5284 25504 5296
rect 25459 5256 25504 5284
rect 25498 5244 25504 5256
rect 25556 5244 25562 5296
rect 30834 5244 30840 5296
rect 30892 5284 30898 5296
rect 31481 5287 31539 5293
rect 31481 5284 31493 5287
rect 30892 5256 31493 5284
rect 30892 5244 30898 5256
rect 31481 5253 31493 5256
rect 31527 5253 31539 5287
rect 33778 5284 33784 5296
rect 33739 5256 33784 5284
rect 31481 5247 31539 5253
rect 33778 5244 33784 5256
rect 33836 5244 33842 5296
rect 25314 5216 25320 5228
rect 25275 5188 25320 5216
rect 25314 5176 25320 5188
rect 25372 5176 25378 5228
rect 27430 5176 27436 5228
rect 27488 5216 27494 5228
rect 27617 5219 27675 5225
rect 27617 5216 27629 5219
rect 27488 5188 27629 5216
rect 27488 5176 27494 5188
rect 27617 5185 27629 5188
rect 27663 5185 27675 5219
rect 27617 5179 27675 5185
rect 28261 5219 28319 5225
rect 28261 5185 28273 5219
rect 28307 5185 28319 5219
rect 28902 5216 28908 5228
rect 28863 5188 28908 5216
rect 28261 5179 28319 5185
rect 24121 5151 24179 5157
rect 24121 5117 24133 5151
rect 24167 5148 24179 5151
rect 24762 5148 24768 5160
rect 24167 5120 24768 5148
rect 24167 5117 24179 5120
rect 24121 5111 24179 5117
rect 24762 5108 24768 5120
rect 24820 5108 24826 5160
rect 26234 5108 26240 5160
rect 26292 5148 26298 5160
rect 26292 5120 26337 5148
rect 26292 5108 26298 5120
rect 26326 5040 26332 5092
rect 26384 5080 26390 5092
rect 28276 5080 28304 5179
rect 28902 5176 28908 5188
rect 28960 5176 28966 5228
rect 28353 5151 28411 5157
rect 28353 5117 28365 5151
rect 28399 5148 28411 5151
rect 29089 5151 29147 5157
rect 29089 5148 29101 5151
rect 28399 5120 29101 5148
rect 28399 5117 28411 5120
rect 28353 5111 28411 5117
rect 29089 5117 29101 5120
rect 29135 5117 29147 5151
rect 30374 5148 30380 5160
rect 30335 5120 30380 5148
rect 29089 5111 29147 5117
rect 30374 5108 30380 5120
rect 30432 5108 30438 5160
rect 31294 5148 31300 5160
rect 31255 5120 31300 5148
rect 31294 5108 31300 5120
rect 31352 5108 31358 5160
rect 31754 5148 31760 5160
rect 31715 5120 31760 5148
rect 31754 5108 31760 5120
rect 31812 5108 31818 5160
rect 33594 5148 33600 5160
rect 33555 5120 33600 5148
rect 33594 5108 33600 5120
rect 33652 5108 33658 5160
rect 34054 5148 34060 5160
rect 34015 5120 34060 5148
rect 34054 5108 34060 5120
rect 34112 5108 34118 5160
rect 28994 5080 29000 5092
rect 26384 5052 29000 5080
rect 26384 5040 26390 5052
rect 28994 5040 29000 5052
rect 29052 5040 29058 5092
rect 23106 4972 23112 5024
rect 23164 5012 23170 5024
rect 23201 5015 23259 5021
rect 23201 5012 23213 5015
rect 23164 4984 23213 5012
rect 23164 4972 23170 4984
rect 23201 4981 23213 4984
rect 23247 4981 23259 5015
rect 23201 4975 23259 4981
rect 24765 5015 24823 5021
rect 24765 4981 24777 5015
rect 24811 5012 24823 5015
rect 25866 5012 25872 5024
rect 24811 4984 25872 5012
rect 24811 4981 24823 4984
rect 24765 4975 24823 4981
rect 25866 4972 25872 4984
rect 25924 4972 25930 5024
rect 36078 5012 36084 5024
rect 36039 4984 36084 5012
rect 36078 4972 36084 4984
rect 36136 4972 36142 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 24765 4811 24823 4817
rect 24765 4777 24777 4811
rect 24811 4808 24823 4811
rect 27890 4808 27896 4820
rect 24811 4780 27896 4808
rect 24811 4777 24823 4780
rect 24765 4771 24823 4777
rect 27890 4768 27896 4780
rect 27948 4768 27954 4820
rect 32769 4811 32827 4817
rect 32769 4777 32781 4811
rect 32815 4808 32827 4811
rect 33594 4808 33600 4820
rect 32815 4780 33600 4808
rect 32815 4777 32827 4780
rect 32769 4771 32827 4777
rect 33594 4768 33600 4780
rect 33652 4768 33658 4820
rect 23477 4743 23535 4749
rect 23477 4709 23489 4743
rect 23523 4740 23535 4743
rect 23934 4740 23940 4752
rect 23523 4712 23940 4740
rect 23523 4709 23535 4712
rect 23477 4703 23535 4709
rect 23934 4700 23940 4712
rect 23992 4700 23998 4752
rect 25409 4743 25467 4749
rect 25409 4709 25421 4743
rect 25455 4740 25467 4743
rect 27246 4740 27252 4752
rect 25455 4712 27252 4740
rect 25455 4709 25467 4712
rect 25409 4703 25467 4709
rect 27246 4700 27252 4712
rect 27304 4700 27310 4752
rect 25866 4672 25872 4684
rect 25827 4644 25872 4672
rect 25866 4632 25872 4644
rect 25924 4632 25930 4684
rect 26418 4672 26424 4684
rect 26379 4644 26424 4672
rect 26418 4632 26424 4644
rect 26476 4632 26482 4684
rect 30742 4672 30748 4684
rect 30703 4644 30748 4672
rect 30742 4632 30748 4644
rect 30800 4632 30806 4684
rect 36078 4672 36084 4684
rect 36039 4644 36084 4672
rect 36078 4632 36084 4644
rect 36136 4632 36142 4684
rect 21450 4564 21456 4616
rect 21508 4604 21514 4616
rect 21545 4607 21603 4613
rect 21545 4604 21557 4607
rect 21508 4576 21557 4604
rect 21508 4564 21514 4576
rect 21545 4573 21557 4576
rect 21591 4573 21603 4607
rect 21545 4567 21603 4573
rect 22554 4564 22560 4616
rect 22612 4604 22618 4616
rect 22649 4607 22707 4613
rect 22649 4604 22661 4607
rect 22612 4576 22661 4604
rect 22612 4564 22618 4576
rect 22649 4573 22661 4576
rect 22695 4573 22707 4607
rect 22649 4567 22707 4573
rect 23937 4607 23995 4613
rect 23937 4573 23949 4607
rect 23983 4604 23995 4607
rect 24118 4604 24124 4616
rect 23983 4576 24124 4604
rect 23983 4573 23995 4576
rect 23937 4567 23995 4573
rect 24118 4564 24124 4576
rect 24176 4564 24182 4616
rect 28534 4604 28540 4616
rect 28495 4576 28540 4604
rect 28534 4564 28540 4576
rect 28592 4564 28598 4616
rect 28994 4604 29000 4616
rect 28955 4576 29000 4604
rect 28994 4564 29000 4576
rect 29052 4564 29058 4616
rect 29825 4607 29883 4613
rect 29825 4573 29837 4607
rect 29871 4604 29883 4607
rect 30285 4607 30343 4613
rect 30285 4604 30297 4607
rect 29871 4576 30297 4604
rect 29871 4573 29883 4576
rect 29825 4567 29883 4573
rect 30285 4573 30297 4576
rect 30331 4573 30343 4607
rect 30285 4567 30343 4573
rect 33413 4607 33471 4613
rect 33413 4573 33425 4607
rect 33459 4604 33471 4607
rect 34514 4604 34520 4616
rect 33459 4576 34520 4604
rect 33459 4573 33471 4576
rect 33413 4567 33471 4573
rect 34514 4564 34520 4576
rect 34572 4564 34578 4616
rect 36722 4604 36728 4616
rect 36683 4576 36728 4604
rect 36722 4564 36728 4576
rect 36780 4564 36786 4616
rect 24029 4539 24087 4545
rect 24029 4505 24041 4539
rect 24075 4536 24087 4539
rect 26053 4539 26111 4545
rect 26053 4536 26065 4539
rect 24075 4508 26065 4536
rect 24075 4505 24087 4508
rect 24029 4499 24087 4505
rect 26053 4505 26065 4508
rect 26099 4505 26111 4539
rect 26053 4499 26111 4505
rect 29089 4539 29147 4545
rect 29089 4505 29101 4539
rect 29135 4536 29147 4539
rect 30469 4539 30527 4545
rect 30469 4536 30481 4539
rect 29135 4508 30481 4536
rect 29135 4505 29147 4508
rect 29089 4499 29147 4505
rect 30469 4505 30481 4508
rect 30515 4505 30527 4539
rect 30469 4499 30527 4505
rect 34146 4496 34152 4548
rect 34204 4536 34210 4548
rect 34241 4539 34299 4545
rect 34241 4536 34253 4539
rect 34204 4508 34253 4536
rect 34204 4496 34210 4508
rect 34241 4505 34253 4508
rect 34287 4505 34299 4539
rect 34241 4499 34299 4505
rect 35897 4539 35955 4545
rect 35897 4505 35909 4539
rect 35943 4536 35955 4539
rect 36633 4539 36691 4545
rect 36633 4536 36645 4539
rect 35943 4508 36645 4536
rect 35943 4505 35955 4508
rect 35897 4499 35955 4505
rect 36633 4505 36645 4508
rect 36679 4505 36691 4539
rect 36633 4499 36691 4505
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 27430 4264 27436 4276
rect 25332 4236 27436 4264
rect 23937 4131 23995 4137
rect 23937 4097 23949 4131
rect 23983 4128 23995 4131
rect 24118 4128 24124 4140
rect 23983 4100 24124 4128
rect 23983 4097 23995 4100
rect 23937 4091 23995 4097
rect 24118 4088 24124 4100
rect 24176 4128 24182 4140
rect 25332 4137 25360 4236
rect 27430 4224 27436 4236
rect 27488 4224 27494 4276
rect 34333 4199 34391 4205
rect 34333 4165 34345 4199
rect 34379 4196 34391 4199
rect 34379 4168 34744 4196
rect 34379 4165 34391 4168
rect 34333 4159 34391 4165
rect 24581 4131 24639 4137
rect 24581 4128 24593 4131
rect 24176 4100 24593 4128
rect 24176 4088 24182 4100
rect 24581 4097 24593 4100
rect 24627 4128 24639 4131
rect 25317 4131 25375 4137
rect 25317 4128 25329 4131
rect 24627 4100 25329 4128
rect 24627 4097 24639 4100
rect 24581 4091 24639 4097
rect 25317 4097 25329 4100
rect 25363 4097 25375 4131
rect 25317 4091 25375 4097
rect 25498 4088 25504 4140
rect 25556 4128 25562 4140
rect 25961 4131 26019 4137
rect 25961 4128 25973 4131
rect 25556 4100 25973 4128
rect 25556 4088 25562 4100
rect 25961 4097 25973 4100
rect 26007 4128 26019 4131
rect 26142 4128 26148 4140
rect 26007 4100 26148 4128
rect 26007 4097 26019 4100
rect 25961 4091 26019 4097
rect 26142 4088 26148 4100
rect 26200 4088 26206 4140
rect 28534 4088 28540 4140
rect 28592 4128 28598 4140
rect 28905 4131 28963 4137
rect 28905 4128 28917 4131
rect 28592 4100 28917 4128
rect 28592 4088 28598 4100
rect 28905 4097 28917 4100
rect 28951 4097 28963 4131
rect 31294 4128 31300 4140
rect 31255 4100 31300 4128
rect 28905 4091 28963 4097
rect 31294 4088 31300 4100
rect 31352 4088 31358 4140
rect 34514 4088 34520 4140
rect 34572 4128 34578 4140
rect 34716 4128 34744 4168
rect 35069 4131 35127 4137
rect 35069 4128 35081 4131
rect 34572 4100 34617 4128
rect 34716 4100 35081 4128
rect 34572 4088 34578 4100
rect 35069 4097 35081 4100
rect 35115 4097 35127 4131
rect 35069 4091 35127 4097
rect 35161 4131 35219 4137
rect 35161 4097 35173 4131
rect 35207 4128 35219 4131
rect 36722 4128 36728 4140
rect 35207 4100 36728 4128
rect 35207 4097 35219 4100
rect 35161 4091 35219 4097
rect 23477 4063 23535 4069
rect 23477 4029 23489 4063
rect 23523 4060 23535 4063
rect 25866 4060 25872 4072
rect 23523 4032 25872 4060
rect 23523 4029 23535 4032
rect 23477 4023 23535 4029
rect 25866 4020 25872 4032
rect 25924 4020 25930 4072
rect 26602 4060 26608 4072
rect 26068 4032 26234 4060
rect 26563 4032 26608 4060
rect 22189 3995 22247 4001
rect 22189 3961 22201 3995
rect 22235 3992 22247 3995
rect 23658 3992 23664 4004
rect 22235 3964 23664 3992
rect 22235 3961 22247 3964
rect 22189 3955 22247 3961
rect 23658 3952 23664 3964
rect 23716 3952 23722 4004
rect 24029 3995 24087 4001
rect 24029 3961 24041 3995
rect 24075 3992 24087 3995
rect 26068 3992 26096 4032
rect 24075 3964 26096 3992
rect 26206 3992 26234 4032
rect 26602 4020 26608 4032
rect 26660 4020 26666 4072
rect 26789 4063 26847 4069
rect 26789 4029 26801 4063
rect 26835 4029 26847 4063
rect 26789 4023 26847 4029
rect 28445 4063 28503 4069
rect 28445 4029 28457 4063
rect 28491 4060 28503 4063
rect 29089 4063 29147 4069
rect 28491 4032 28948 4060
rect 28491 4029 28503 4032
rect 28445 4023 28503 4029
rect 26804 3992 26832 4023
rect 28920 4004 28948 4032
rect 29089 4029 29101 4063
rect 29135 4029 29147 4063
rect 29730 4060 29736 4072
rect 29691 4032 29736 4060
rect 29089 4023 29147 4029
rect 26206 3964 26832 3992
rect 24075 3961 24087 3964
rect 24029 3955 24087 3961
rect 28902 3952 28908 4004
rect 28960 3952 28966 4004
rect 19889 3927 19947 3933
rect 19889 3893 19901 3927
rect 19935 3924 19947 3927
rect 19978 3924 19984 3936
rect 19935 3896 19984 3924
rect 19935 3893 19947 3896
rect 19889 3887 19947 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 20717 3927 20775 3933
rect 20717 3924 20729 3927
rect 20680 3896 20729 3924
rect 20680 3884 20686 3896
rect 20717 3893 20729 3896
rect 20763 3893 20775 3927
rect 20717 3887 20775 3893
rect 21545 3927 21603 3933
rect 21545 3893 21557 3927
rect 21591 3924 21603 3927
rect 22002 3924 22008 3936
rect 21591 3896 22008 3924
rect 21591 3893 21603 3896
rect 21545 3887 21603 3893
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 22833 3927 22891 3933
rect 22833 3893 22845 3927
rect 22879 3924 22891 3927
rect 24486 3924 24492 3936
rect 22879 3896 24492 3924
rect 22879 3893 22891 3896
rect 22833 3887 22891 3893
rect 24486 3884 24492 3896
rect 24544 3884 24550 3936
rect 24670 3924 24676 3936
rect 24631 3896 24676 3924
rect 24670 3884 24676 3896
rect 24728 3884 24734 3936
rect 25406 3924 25412 3936
rect 25367 3896 25412 3924
rect 25406 3884 25412 3896
rect 25464 3884 25470 3936
rect 26050 3924 26056 3936
rect 26011 3896 26056 3924
rect 26050 3884 26056 3896
rect 26108 3884 26114 3936
rect 26142 3884 26148 3936
rect 26200 3924 26206 3936
rect 26326 3924 26332 3936
rect 26200 3896 26332 3924
rect 26200 3884 26206 3896
rect 26326 3884 26332 3896
rect 26384 3884 26390 3936
rect 26510 3884 26516 3936
rect 26568 3924 26574 3936
rect 29104 3924 29132 4023
rect 29730 4020 29736 4032
rect 29788 4020 29794 4072
rect 33042 4060 33048 4072
rect 33003 4032 33048 4060
rect 33042 4020 33048 4032
rect 33100 4020 33106 4072
rect 35176 4060 35204 4091
rect 36722 4088 36728 4100
rect 36780 4088 36786 4140
rect 34256 4032 35204 4060
rect 30466 3952 30472 4004
rect 30524 3992 30530 4004
rect 34256 3992 34284 4032
rect 30524 3964 34284 3992
rect 30524 3952 30530 3964
rect 37182 3952 37188 4004
rect 37240 3992 37246 4004
rect 37921 3995 37979 4001
rect 37921 3992 37933 3995
rect 37240 3964 37933 3992
rect 37240 3952 37246 3964
rect 37921 3961 37933 3964
rect 37967 3961 37979 3995
rect 37921 3955 37979 3961
rect 26568 3896 29132 3924
rect 26568 3884 26574 3896
rect 31478 3884 31484 3936
rect 31536 3924 31542 3936
rect 31941 3927 31999 3933
rect 31941 3924 31953 3927
rect 31536 3896 31953 3924
rect 31536 3884 31542 3896
rect 31941 3893 31953 3896
rect 31987 3893 31999 3927
rect 31941 3887 31999 3893
rect 33410 3884 33416 3936
rect 33468 3924 33474 3936
rect 35621 3927 35679 3933
rect 35621 3924 35633 3927
rect 33468 3896 35633 3924
rect 33468 3884 33474 3896
rect 35621 3893 35633 3896
rect 35667 3893 35679 3927
rect 35621 3887 35679 3893
rect 35710 3884 35716 3936
rect 35768 3924 35774 3936
rect 36265 3927 36323 3933
rect 36265 3924 36277 3927
rect 35768 3896 36277 3924
rect 35768 3884 35774 3896
rect 36265 3893 36277 3896
rect 36311 3893 36323 3927
rect 37274 3924 37280 3936
rect 37235 3896 37280 3924
rect 36265 3887 36323 3893
rect 37274 3884 37280 3896
rect 37332 3884 37338 3936
rect 38562 3884 38568 3936
rect 38620 3924 38626 3936
rect 38657 3927 38715 3933
rect 38657 3924 38669 3927
rect 38620 3896 38669 3924
rect 38620 3884 38626 3896
rect 38657 3893 38669 3896
rect 38703 3893 38715 3927
rect 38657 3887 38715 3893
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 22830 3680 22836 3732
rect 22888 3720 22894 3732
rect 26602 3720 26608 3732
rect 22888 3692 26608 3720
rect 22888 3680 22894 3692
rect 26602 3680 26608 3692
rect 26660 3680 26666 3732
rect 30834 3720 30840 3732
rect 30795 3692 30840 3720
rect 30834 3680 30840 3692
rect 30892 3680 30898 3732
rect 36078 3680 36084 3732
rect 36136 3720 36142 3732
rect 37829 3723 37887 3729
rect 37829 3720 37841 3723
rect 36136 3692 37841 3720
rect 36136 3680 36142 3692
rect 37829 3689 37841 3692
rect 37875 3689 37887 3723
rect 37829 3683 37887 3689
rect 21085 3655 21143 3661
rect 21085 3621 21097 3655
rect 21131 3652 21143 3655
rect 22278 3652 22284 3664
rect 21131 3624 22284 3652
rect 21131 3621 21143 3624
rect 21085 3615 21143 3621
rect 22278 3612 22284 3624
rect 22336 3612 22342 3664
rect 24118 3652 24124 3664
rect 22940 3624 24124 3652
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 9401 3519 9459 3525
rect 9401 3516 9413 3519
rect 9364 3488 9413 3516
rect 9364 3476 9370 3488
rect 9401 3485 9413 3488
rect 9447 3485 9459 3519
rect 9401 3479 9459 3485
rect 10778 3476 10784 3528
rect 10836 3516 10842 3528
rect 10873 3519 10931 3525
rect 10873 3516 10885 3519
rect 10836 3488 10885 3516
rect 10836 3476 10842 3488
rect 10873 3485 10885 3488
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 12529 3519 12587 3525
rect 12529 3516 12541 3519
rect 12492 3488 12541 3516
rect 12492 3476 12498 3488
rect 12529 3485 12541 3488
rect 12575 3485 12587 3519
rect 12529 3479 12587 3485
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 13633 3519 13691 3525
rect 13633 3516 13645 3519
rect 13596 3488 13645 3516
rect 13596 3476 13602 3488
rect 13633 3485 13645 3488
rect 13679 3485 13691 3519
rect 13633 3479 13691 3485
rect 14642 3476 14648 3528
rect 14700 3516 14706 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14700 3488 14749 3516
rect 14700 3476 14706 3488
rect 14737 3485 14749 3488
rect 14783 3485 14795 3519
rect 14737 3479 14795 3485
rect 15470 3476 15476 3528
rect 15528 3516 15534 3528
rect 15565 3519 15623 3525
rect 15565 3516 15577 3519
rect 15528 3488 15577 3516
rect 15528 3476 15534 3488
rect 15565 3485 15577 3488
rect 15611 3485 15623 3519
rect 15565 3479 15623 3485
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 16632 3488 16681 3516
rect 16632 3476 16638 3488
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 17310 3476 17316 3528
rect 17368 3516 17374 3528
rect 17405 3519 17463 3525
rect 17405 3516 17417 3519
rect 17368 3488 17417 3516
rect 17368 3476 17374 3488
rect 17405 3485 17417 3488
rect 17451 3485 17463 3519
rect 17405 3479 17463 3485
rect 18138 3476 18144 3528
rect 18196 3516 18202 3528
rect 18233 3519 18291 3525
rect 18233 3516 18245 3519
rect 18196 3488 18245 3516
rect 18196 3476 18202 3488
rect 18233 3485 18245 3488
rect 18279 3485 18291 3519
rect 18966 3516 18972 3528
rect 18927 3488 18972 3516
rect 18233 3479 18291 3485
rect 18966 3476 18972 3488
rect 19024 3476 19030 3528
rect 19797 3519 19855 3525
rect 19797 3485 19809 3519
rect 19843 3516 19855 3519
rect 20346 3516 20352 3528
rect 19843 3488 20352 3516
rect 19843 3485 19855 3488
rect 19797 3479 19855 3485
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 20441 3519 20499 3525
rect 20441 3485 20453 3519
rect 20487 3516 20499 3519
rect 20898 3516 20904 3528
rect 20487 3488 20904 3516
rect 20487 3485 20499 3488
rect 20441 3479 20499 3485
rect 20898 3476 20904 3488
rect 20956 3476 20962 3528
rect 21729 3519 21787 3525
rect 21729 3485 21741 3519
rect 21775 3485 21787 3519
rect 21729 3479 21787 3485
rect 21744 3380 21772 3479
rect 22186 3476 22192 3528
rect 22244 3516 22250 3528
rect 22940 3525 22968 3624
rect 24118 3612 24124 3624
rect 24176 3612 24182 3664
rect 24486 3612 24492 3664
rect 24544 3652 24550 3664
rect 25314 3652 25320 3664
rect 24544 3624 25320 3652
rect 24544 3612 24550 3624
rect 25314 3612 25320 3624
rect 25372 3612 25378 3664
rect 25406 3612 25412 3664
rect 25464 3652 25470 3664
rect 25464 3624 26234 3652
rect 25464 3612 25470 3624
rect 23017 3587 23075 3593
rect 23017 3553 23029 3587
rect 23063 3584 23075 3587
rect 26053 3587 26111 3593
rect 26053 3584 26065 3587
rect 23063 3556 26065 3584
rect 23063 3553 23075 3556
rect 23017 3547 23075 3553
rect 26053 3553 26065 3556
rect 26099 3553 26111 3587
rect 26206 3584 26234 3624
rect 28350 3612 28356 3664
rect 28408 3652 28414 3664
rect 28408 3624 28764 3652
rect 28408 3612 28414 3624
rect 28736 3593 28764 3624
rect 36538 3612 36544 3664
rect 36596 3652 36602 3664
rect 37185 3655 37243 3661
rect 37185 3652 37197 3655
rect 36596 3624 37197 3652
rect 36596 3612 36602 3624
rect 37185 3621 37197 3624
rect 37231 3621 37243 3655
rect 37185 3615 37243 3621
rect 39942 3612 39948 3664
rect 40000 3652 40006 3664
rect 40865 3655 40923 3661
rect 40865 3652 40877 3655
rect 40000 3624 40877 3652
rect 40000 3612 40006 3624
rect 40865 3621 40877 3624
rect 40911 3621 40923 3655
rect 40865 3615 40923 3621
rect 28445 3587 28503 3593
rect 28445 3584 28457 3587
rect 26206 3556 28457 3584
rect 26053 3547 26111 3553
rect 28445 3553 28457 3556
rect 28491 3553 28503 3587
rect 28445 3547 28503 3553
rect 28721 3587 28779 3593
rect 28721 3553 28733 3587
rect 28767 3553 28779 3587
rect 28721 3547 28779 3553
rect 28994 3544 29000 3596
rect 29052 3584 29058 3596
rect 31478 3584 31484 3596
rect 29052 3556 30788 3584
rect 31439 3556 31484 3584
rect 29052 3544 29058 3556
rect 22281 3519 22339 3525
rect 22281 3516 22293 3519
rect 22244 3488 22293 3516
rect 22244 3476 22250 3488
rect 22281 3485 22293 3488
rect 22327 3516 22339 3519
rect 22925 3519 22983 3525
rect 22925 3516 22937 3519
rect 22327 3488 22937 3516
rect 22327 3485 22339 3488
rect 22281 3479 22339 3485
rect 22925 3485 22937 3488
rect 22971 3485 22983 3519
rect 23566 3516 23572 3528
rect 23527 3488 23572 3516
rect 22925 3479 22983 3485
rect 23566 3476 23572 3488
rect 23624 3476 23630 3528
rect 25866 3516 25872 3528
rect 25827 3488 25872 3516
rect 25866 3476 25872 3488
rect 25924 3476 25930 3528
rect 27246 3476 27252 3528
rect 27304 3516 27310 3528
rect 30760 3525 30788 3556
rect 31478 3544 31484 3556
rect 31536 3544 31542 3596
rect 31938 3584 31944 3596
rect 31899 3556 31944 3584
rect 31938 3544 31944 3556
rect 31996 3544 32002 3596
rect 34422 3584 34428 3596
rect 34383 3556 34428 3584
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 36081 3587 36139 3593
rect 36081 3553 36093 3587
rect 36127 3584 36139 3587
rect 37274 3584 37280 3596
rect 36127 3556 37280 3584
rect 36127 3553 36139 3556
rect 36081 3547 36139 3553
rect 37274 3544 37280 3556
rect 37332 3544 37338 3596
rect 37550 3544 37556 3596
rect 37608 3584 37614 3596
rect 39117 3587 39175 3593
rect 39117 3584 39129 3587
rect 37608 3556 39129 3584
rect 37608 3544 37614 3556
rect 39117 3553 39129 3556
rect 39163 3553 39175 3587
rect 39117 3547 39175 3553
rect 40770 3544 40776 3596
rect 40828 3584 40834 3596
rect 41509 3587 41567 3593
rect 41509 3584 41521 3587
rect 40828 3556 41521 3584
rect 40828 3544 40834 3556
rect 41509 3553 41521 3556
rect 41555 3553 41567 3587
rect 41509 3547 41567 3553
rect 28261 3519 28319 3525
rect 28261 3516 28273 3519
rect 27304 3488 28273 3516
rect 27304 3476 27310 3488
rect 28261 3485 28273 3488
rect 28307 3485 28319 3519
rect 28261 3479 28319 3485
rect 30745 3519 30803 3525
rect 30745 3485 30757 3519
rect 30791 3485 30803 3519
rect 36722 3516 36728 3528
rect 36683 3488 36728 3516
rect 30745 3479 30803 3485
rect 36722 3476 36728 3488
rect 36780 3476 36786 3528
rect 36814 3476 36820 3528
rect 36872 3516 36878 3528
rect 38473 3519 38531 3525
rect 38473 3516 38485 3519
rect 36872 3488 38485 3516
rect 36872 3476 36878 3488
rect 38473 3485 38485 3488
rect 38519 3485 38531 3519
rect 38473 3479 38531 3485
rect 39390 3476 39396 3528
rect 39448 3516 39454 3528
rect 40221 3519 40279 3525
rect 40221 3516 40233 3519
rect 39448 3488 40233 3516
rect 39448 3476 39454 3488
rect 40221 3485 40233 3488
rect 40267 3485 40279 3519
rect 40221 3479 40279 3485
rect 41322 3476 41328 3528
rect 41380 3516 41386 3528
rect 42153 3519 42211 3525
rect 42153 3516 42165 3519
rect 41380 3488 42165 3516
rect 41380 3476 41386 3488
rect 42153 3485 42165 3488
rect 42199 3485 42211 3519
rect 42153 3479 42211 3485
rect 42426 3476 42432 3528
rect 42484 3516 42490 3528
rect 42797 3519 42855 3525
rect 42797 3516 42809 3519
rect 42484 3488 42809 3516
rect 42484 3476 42490 3488
rect 42797 3485 42809 3488
rect 42843 3485 42855 3519
rect 42797 3479 42855 3485
rect 43254 3476 43260 3528
rect 43312 3516 43318 3528
rect 43441 3519 43499 3525
rect 43441 3516 43453 3519
rect 43312 3488 43453 3516
rect 43312 3476 43318 3488
rect 43441 3485 43453 3488
rect 43487 3485 43499 3519
rect 43441 3479 43499 3485
rect 44082 3476 44088 3528
rect 44140 3516 44146 3528
rect 44177 3519 44235 3525
rect 44177 3516 44189 3519
rect 44140 3488 44189 3516
rect 44140 3476 44146 3488
rect 44177 3485 44189 3488
rect 44223 3485 44235 3519
rect 44177 3479 44235 3485
rect 46014 3476 46020 3528
rect 46072 3516 46078 3528
rect 46201 3519 46259 3525
rect 46201 3516 46213 3519
rect 46072 3488 46213 3516
rect 46072 3476 46078 3488
rect 46201 3485 46213 3488
rect 46247 3485 46259 3519
rect 46201 3479 46259 3485
rect 46566 3476 46572 3528
rect 46624 3516 46630 3528
rect 46845 3519 46903 3525
rect 46845 3516 46857 3519
rect 46624 3488 46857 3516
rect 46624 3476 46630 3488
rect 46845 3485 46857 3488
rect 46891 3485 46903 3519
rect 46845 3479 46903 3485
rect 48222 3476 48228 3528
rect 48280 3516 48286 3528
rect 48317 3519 48375 3525
rect 48317 3516 48329 3519
rect 48280 3488 48329 3516
rect 48280 3476 48286 3488
rect 48317 3485 48329 3488
rect 48363 3485 48375 3519
rect 48317 3479 48375 3485
rect 49326 3476 49332 3528
rect 49384 3516 49390 3528
rect 49421 3519 49479 3525
rect 49421 3516 49433 3519
rect 49384 3488 49433 3516
rect 49384 3476 49390 3488
rect 49421 3485 49433 3488
rect 49467 3485 49479 3519
rect 49421 3479 49479 3485
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50249 3519 50307 3525
rect 50249 3516 50261 3519
rect 50212 3488 50261 3516
rect 50212 3476 50218 3488
rect 50249 3485 50261 3488
rect 50295 3485 50307 3519
rect 50249 3479 50307 3485
rect 52086 3476 52092 3528
rect 52144 3516 52150 3528
rect 52181 3519 52239 3525
rect 52181 3516 52193 3519
rect 52144 3488 52193 3516
rect 52144 3476 52150 3488
rect 52181 3485 52193 3488
rect 52227 3485 52239 3519
rect 52181 3479 52239 3485
rect 22373 3451 22431 3457
rect 22373 3417 22385 3451
rect 22419 3448 22431 3451
rect 23753 3451 23811 3457
rect 23753 3448 23765 3451
rect 22419 3420 23765 3448
rect 22419 3417 22431 3420
rect 22373 3411 22431 3417
rect 23753 3417 23765 3420
rect 23799 3417 23811 3451
rect 23753 3411 23811 3417
rect 25409 3451 25467 3457
rect 25409 3417 25421 3451
rect 25455 3448 25467 3451
rect 25455 3420 26648 3448
rect 25455 3417 25467 3420
rect 25409 3411 25467 3417
rect 24302 3380 24308 3392
rect 21744 3352 24308 3380
rect 24302 3340 24308 3352
rect 24360 3340 24366 3392
rect 26050 3340 26056 3392
rect 26108 3380 26114 3392
rect 26510 3380 26516 3392
rect 26108 3352 26516 3380
rect 26108 3340 26114 3352
rect 26510 3340 26516 3352
rect 26568 3340 26574 3392
rect 26620 3380 26648 3420
rect 26694 3408 26700 3460
rect 26752 3448 26758 3460
rect 27709 3451 27767 3457
rect 27709 3448 27721 3451
rect 26752 3420 27721 3448
rect 26752 3408 26758 3420
rect 27709 3417 27721 3420
rect 27755 3417 27767 3451
rect 27709 3411 27767 3417
rect 27798 3408 27804 3460
rect 27856 3448 27862 3460
rect 29178 3448 29184 3460
rect 27856 3420 29184 3448
rect 27856 3408 27862 3420
rect 29178 3408 29184 3420
rect 29236 3408 29242 3460
rect 30650 3408 30656 3460
rect 30708 3448 30714 3460
rect 31665 3451 31723 3457
rect 31665 3448 31677 3451
rect 30708 3420 31677 3448
rect 30708 3408 30714 3420
rect 31665 3417 31677 3420
rect 31711 3417 31723 3451
rect 31665 3411 31723 3417
rect 35897 3451 35955 3457
rect 35897 3417 35909 3451
rect 35943 3448 35955 3451
rect 37458 3448 37464 3460
rect 35943 3420 37464 3448
rect 35943 3417 35955 3420
rect 35897 3411 35955 3417
rect 37458 3408 37464 3420
rect 37516 3408 37522 3460
rect 26970 3380 26976 3392
rect 26620 3352 26976 3380
rect 26970 3340 26976 3352
rect 27028 3340 27034 3392
rect 33226 3340 33232 3392
rect 33284 3380 33290 3392
rect 36633 3383 36691 3389
rect 36633 3380 36645 3383
rect 33284 3352 36645 3380
rect 33284 3340 33290 3352
rect 36633 3349 36645 3352
rect 36679 3349 36691 3383
rect 36633 3343 36691 3349
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 24670 3136 24676 3188
rect 24728 3176 24734 3188
rect 30650 3176 30656 3188
rect 24728 3148 26234 3176
rect 30611 3148 30656 3176
rect 24728 3136 24734 3148
rect 23385 3111 23443 3117
rect 23385 3077 23397 3111
rect 23431 3108 23443 3111
rect 25777 3111 25835 3117
rect 25777 3108 25789 3111
rect 23431 3080 25789 3108
rect 23431 3077 23443 3080
rect 23385 3071 23443 3077
rect 25777 3077 25789 3080
rect 25823 3077 25835 3111
rect 26206 3108 26234 3148
rect 30650 3136 30656 3148
rect 30708 3136 30714 3188
rect 28077 3111 28135 3117
rect 28077 3108 28089 3111
rect 26206 3080 28089 3108
rect 25777 3071 25835 3077
rect 28077 3077 28089 3080
rect 28123 3077 28135 3111
rect 33226 3108 33232 3120
rect 33187 3080 33232 3108
rect 28077 3071 28135 3077
rect 33226 3068 33232 3080
rect 33284 3068 33290 3120
rect 35529 3111 35587 3117
rect 35529 3077 35541 3111
rect 35575 3108 35587 3111
rect 37369 3111 37427 3117
rect 37369 3108 37381 3111
rect 35575 3080 37381 3108
rect 35575 3077 35587 3080
rect 35529 3071 35587 3077
rect 37369 3077 37381 3080
rect 37415 3077 37427 3111
rect 37369 3071 37427 3077
rect 20901 3043 20959 3049
rect 20901 3009 20913 3043
rect 20947 3040 20959 3043
rect 20947 3012 22140 3040
rect 20947 3009 20959 3012
rect 20901 3003 20959 3009
rect 16209 2975 16267 2981
rect 16209 2941 16221 2975
rect 16255 2972 16267 2975
rect 16850 2972 16856 2984
rect 16255 2944 16856 2972
rect 16255 2941 16267 2944
rect 16209 2935 16267 2941
rect 16850 2932 16856 2944
rect 16908 2932 16914 2984
rect 19613 2975 19671 2981
rect 19613 2941 19625 2975
rect 19659 2972 19671 2975
rect 21174 2972 21180 2984
rect 19659 2944 21180 2972
rect 19659 2941 19671 2944
rect 19613 2935 19671 2941
rect 21174 2932 21180 2944
rect 21232 2932 21238 2984
rect 22112 2972 22140 3012
rect 22186 3000 22192 3052
rect 22244 3040 22250 3052
rect 22830 3040 22836 3052
rect 22244 3012 22289 3040
rect 22791 3012 22836 3040
rect 22244 3000 22250 3012
rect 22830 3000 22836 3012
rect 22888 3000 22894 3052
rect 23477 3043 23535 3049
rect 23477 3009 23489 3043
rect 23523 3040 23535 3043
rect 24210 3040 24216 3052
rect 23523 3012 24216 3040
rect 23523 3009 23535 3012
rect 23477 3003 23535 3009
rect 24210 3000 24216 3012
rect 24268 3040 24274 3052
rect 24581 3043 24639 3049
rect 24581 3040 24593 3043
rect 24268 3012 24593 3040
rect 24268 3000 24274 3012
rect 24581 3009 24593 3012
rect 24627 3040 24639 3043
rect 25498 3040 25504 3052
rect 24627 3012 25504 3040
rect 24627 3009 24639 3012
rect 24581 3003 24639 3009
rect 25498 3000 25504 3012
rect 25556 3000 25562 3052
rect 27614 3040 27620 3052
rect 27356 3012 27620 3040
rect 23382 2972 23388 2984
rect 22112 2944 23388 2972
rect 23382 2932 23388 2944
rect 23440 2932 23446 2984
rect 24670 2972 24676 2984
rect 24631 2944 24676 2972
rect 24670 2932 24676 2944
rect 24728 2932 24734 2984
rect 25590 2972 25596 2984
rect 25551 2944 25596 2972
rect 25590 2932 25596 2944
rect 25648 2932 25654 2984
rect 20257 2907 20315 2913
rect 20257 2873 20269 2907
rect 20303 2904 20315 2907
rect 21726 2904 21732 2916
rect 20303 2876 21732 2904
rect 20303 2873 20315 2876
rect 20257 2867 20315 2873
rect 21726 2864 21732 2876
rect 21784 2864 21790 2916
rect 22097 2907 22155 2913
rect 22097 2873 22109 2907
rect 22143 2904 22155 2907
rect 24026 2904 24032 2916
rect 22143 2876 24032 2904
rect 22143 2873 22155 2876
rect 22097 2867 22155 2873
rect 24026 2864 24032 2876
rect 24084 2864 24090 2916
rect 24121 2907 24179 2913
rect 24121 2873 24133 2907
rect 24167 2904 24179 2907
rect 27356 2904 27384 3012
rect 27614 3000 27620 3012
rect 27672 3000 27678 3052
rect 27890 3040 27896 3052
rect 27851 3012 27896 3040
rect 27890 3000 27896 3012
rect 27948 3000 27954 3052
rect 30466 3000 30472 3052
rect 30524 3040 30530 3052
rect 30561 3043 30619 3049
rect 30561 3040 30573 3043
rect 30524 3012 30573 3040
rect 30524 3000 30530 3012
rect 30561 3009 30573 3012
rect 30607 3009 30619 3043
rect 30561 3003 30619 3009
rect 31386 3000 31392 3052
rect 31444 3040 31450 3052
rect 31754 3040 31760 3052
rect 31444 3012 31760 3040
rect 31444 3000 31450 3012
rect 31754 3000 31760 3012
rect 31812 3000 31818 3052
rect 33410 3000 33416 3052
rect 33468 3040 33474 3052
rect 33468 3012 33513 3040
rect 33468 3000 33474 3012
rect 35710 3000 35716 3052
rect 35768 3040 35774 3052
rect 35768 3012 35813 3040
rect 35768 3000 35774 3012
rect 36722 3000 36728 3052
rect 36780 3040 36786 3052
rect 37277 3043 37335 3049
rect 37277 3040 37289 3043
rect 36780 3012 37289 3040
rect 36780 3000 36786 3012
rect 37277 3009 37289 3012
rect 37323 3009 37335 3043
rect 37277 3003 37335 3009
rect 38010 3000 38016 3052
rect 38068 3040 38074 3052
rect 39853 3043 39911 3049
rect 39853 3040 39865 3043
rect 38068 3012 39865 3040
rect 38068 3000 38074 3012
rect 39853 3009 39865 3012
rect 39899 3009 39911 3043
rect 39853 3003 39911 3009
rect 40218 3000 40224 3052
rect 40276 3040 40282 3052
rect 41785 3043 41843 3049
rect 41785 3040 41797 3043
rect 40276 3012 41797 3040
rect 40276 3000 40282 3012
rect 41785 3009 41797 3012
rect 41831 3009 41843 3043
rect 41785 3003 41843 3009
rect 27433 2975 27491 2981
rect 27433 2941 27445 2975
rect 27479 2941 27491 2975
rect 28626 2972 28632 2984
rect 28587 2944 28632 2972
rect 27433 2935 27491 2941
rect 24167 2876 27384 2904
rect 24167 2873 24179 2876
rect 24121 2867 24179 2873
rect 7650 2796 7656 2848
rect 7708 2836 7714 2848
rect 7745 2839 7803 2845
rect 7745 2836 7757 2839
rect 7708 2808 7757 2836
rect 7708 2796 7714 2808
rect 7745 2805 7757 2808
rect 7791 2805 7803 2839
rect 7745 2799 7803 2805
rect 8570 2796 8576 2848
rect 8628 2836 8634 2848
rect 8665 2839 8723 2845
rect 8665 2836 8677 2839
rect 8628 2808 8677 2836
rect 8628 2796 8634 2808
rect 8665 2805 8677 2808
rect 8711 2805 8723 2839
rect 8665 2799 8723 2805
rect 9585 2839 9643 2845
rect 9585 2805 9597 2839
rect 9631 2836 9643 2839
rect 9950 2836 9956 2848
rect 9631 2808 9956 2836
rect 9631 2805 9643 2808
rect 9585 2799 9643 2805
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 10229 2839 10287 2845
rect 10229 2805 10241 2839
rect 10275 2836 10287 2839
rect 10502 2836 10508 2848
rect 10275 2808 10508 2836
rect 10275 2805 10287 2808
rect 10229 2799 10287 2805
rect 10502 2796 10508 2808
rect 10560 2796 10566 2848
rect 10873 2839 10931 2845
rect 10873 2805 10885 2839
rect 10919 2836 10931 2839
rect 11054 2836 11060 2848
rect 10919 2808 11060 2836
rect 10919 2805 10931 2808
rect 10873 2799 10931 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2836 11575 2839
rect 11606 2836 11612 2848
rect 11563 2808 11612 2836
rect 11563 2805 11575 2808
rect 11517 2799 11575 2805
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 12158 2836 12164 2848
rect 12119 2808 12164 2836
rect 12158 2796 12164 2808
rect 12216 2796 12222 2848
rect 12805 2839 12863 2845
rect 12805 2805 12817 2839
rect 12851 2836 12863 2839
rect 12986 2836 12992 2848
rect 12851 2808 12992 2836
rect 12851 2805 12863 2808
rect 12805 2799 12863 2805
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 13633 2839 13691 2845
rect 13633 2805 13645 2839
rect 13679 2836 13691 2839
rect 13814 2836 13820 2848
rect 13679 2808 13820 2836
rect 13679 2805 13691 2808
rect 13633 2799 13691 2805
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 14277 2839 14335 2845
rect 14277 2805 14289 2839
rect 14323 2836 14335 2839
rect 14366 2836 14372 2848
rect 14323 2808 14372 2836
rect 14323 2805 14335 2808
rect 14277 2799 14335 2805
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 14921 2839 14979 2845
rect 14921 2805 14933 2839
rect 14967 2836 14979 2839
rect 15194 2836 15200 2848
rect 14967 2808 15200 2836
rect 14967 2805 14979 2808
rect 14921 2799 14979 2805
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 15565 2839 15623 2845
rect 15565 2805 15577 2839
rect 15611 2836 15623 2839
rect 16022 2836 16028 2848
rect 15611 2808 16028 2836
rect 15611 2805 15623 2808
rect 15565 2799 15623 2805
rect 16022 2796 16028 2808
rect 16080 2796 16086 2848
rect 16853 2839 16911 2845
rect 16853 2805 16865 2839
rect 16899 2836 16911 2839
rect 17126 2836 17132 2848
rect 16899 2808 17132 2836
rect 16899 2805 16911 2808
rect 16853 2799 16911 2805
rect 17126 2796 17132 2808
rect 17184 2796 17190 2848
rect 17497 2839 17555 2845
rect 17497 2805 17509 2839
rect 17543 2836 17555 2839
rect 17862 2836 17868 2848
rect 17543 2808 17868 2836
rect 17543 2805 17555 2808
rect 17497 2799 17555 2805
rect 17862 2796 17868 2808
rect 17920 2796 17926 2848
rect 18141 2839 18199 2845
rect 18141 2805 18153 2839
rect 18187 2836 18199 2839
rect 18690 2836 18696 2848
rect 18187 2808 18696 2836
rect 18187 2805 18199 2808
rect 18141 2799 18199 2805
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 18785 2839 18843 2845
rect 18785 2805 18797 2839
rect 18831 2836 18843 2839
rect 19426 2836 19432 2848
rect 18831 2808 19432 2836
rect 18831 2805 18843 2808
rect 18785 2799 18843 2805
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 21545 2839 21603 2845
rect 21545 2805 21557 2839
rect 21591 2836 21603 2839
rect 25498 2836 25504 2848
rect 21591 2808 25504 2836
rect 21591 2805 21603 2808
rect 21545 2799 21603 2805
rect 25498 2796 25504 2808
rect 25556 2796 25562 2848
rect 27448 2836 27476 2935
rect 28626 2932 28632 2944
rect 28684 2932 28690 2984
rect 32214 2972 32220 2984
rect 32175 2944 32220 2972
rect 32214 2932 32220 2944
rect 32272 2932 32278 2984
rect 33873 2975 33931 2981
rect 33873 2941 33885 2975
rect 33919 2941 33931 2975
rect 33873 2935 33931 2941
rect 33318 2864 33324 2916
rect 33376 2904 33382 2916
rect 33888 2904 33916 2935
rect 35342 2932 35348 2984
rect 35400 2972 35406 2984
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 35400 2944 37933 2972
rect 35400 2932 35406 2944
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 37921 2935 37979 2941
rect 39666 2932 39672 2984
rect 39724 2972 39730 2984
rect 41141 2975 41199 2981
rect 41141 2972 41153 2975
rect 39724 2944 41153 2972
rect 39724 2932 39730 2944
rect 41141 2941 41153 2944
rect 41187 2941 41199 2975
rect 41141 2935 41199 2941
rect 45462 2932 45468 2984
rect 45520 2972 45526 2984
rect 46477 2975 46535 2981
rect 46477 2972 46489 2975
rect 45520 2944 46489 2972
rect 45520 2932 45526 2944
rect 46477 2941 46489 2944
rect 46523 2941 46535 2975
rect 46477 2935 46535 2941
rect 46842 2932 46848 2984
rect 46900 2972 46906 2984
rect 47765 2975 47823 2981
rect 47765 2972 47777 2975
rect 46900 2944 47777 2972
rect 46900 2932 46906 2944
rect 47765 2941 47777 2944
rect 47811 2941 47823 2975
rect 47765 2935 47823 2941
rect 33376 2876 33916 2904
rect 33376 2864 33382 2876
rect 35802 2864 35808 2916
rect 35860 2904 35866 2916
rect 38565 2907 38623 2913
rect 38565 2904 38577 2907
rect 35860 2876 38577 2904
rect 35860 2864 35866 2876
rect 38565 2873 38577 2876
rect 38611 2873 38623 2907
rect 38565 2867 38623 2873
rect 38838 2864 38844 2916
rect 38896 2904 38902 2916
rect 40497 2907 40555 2913
rect 40497 2904 40509 2907
rect 38896 2876 40509 2904
rect 38896 2864 38902 2876
rect 40497 2873 40509 2876
rect 40543 2873 40555 2907
rect 40497 2867 40555 2873
rect 41046 2864 41052 2916
rect 41104 2904 41110 2916
rect 42429 2907 42487 2913
rect 42429 2904 42441 2907
rect 41104 2876 42441 2904
rect 41104 2864 41110 2876
rect 42429 2873 42441 2876
rect 42475 2873 42487 2907
rect 42429 2867 42487 2873
rect 42978 2864 42984 2916
rect 43036 2904 43042 2916
rect 43901 2907 43959 2913
rect 43901 2904 43913 2907
rect 43036 2876 43913 2904
rect 43036 2864 43042 2876
rect 43901 2873 43913 2876
rect 43947 2873 43959 2907
rect 43901 2867 43959 2873
rect 44358 2864 44364 2916
rect 44416 2904 44422 2916
rect 45189 2907 45247 2913
rect 45189 2904 45201 2907
rect 44416 2876 45201 2904
rect 44416 2864 44422 2876
rect 45189 2873 45201 2876
rect 45235 2873 45247 2907
rect 45189 2867 45247 2873
rect 47670 2864 47676 2916
rect 47728 2904 47734 2916
rect 48409 2907 48467 2913
rect 48409 2904 48421 2907
rect 47728 2876 48421 2904
rect 47728 2864 47734 2876
rect 48409 2873 48421 2876
rect 48455 2873 48467 2907
rect 48409 2867 48467 2873
rect 49050 2864 49056 2916
rect 49108 2904 49114 2916
rect 49881 2907 49939 2913
rect 49881 2904 49893 2907
rect 49108 2876 49893 2904
rect 49108 2864 49114 2876
rect 49881 2873 49893 2876
rect 49927 2873 49939 2907
rect 49881 2867 49939 2873
rect 50982 2864 50988 2916
rect 51040 2904 51046 2916
rect 51813 2907 51871 2913
rect 51813 2904 51825 2907
rect 51040 2876 51825 2904
rect 51040 2864 51046 2876
rect 51813 2873 51825 2876
rect 51859 2873 51871 2907
rect 51813 2867 51871 2873
rect 52362 2864 52368 2916
rect 52420 2904 52426 2916
rect 53101 2907 53159 2913
rect 53101 2904 53113 2907
rect 52420 2876 53113 2904
rect 52420 2864 52426 2876
rect 53101 2873 53113 2876
rect 53147 2873 53159 2907
rect 53101 2867 53159 2873
rect 29178 2836 29184 2848
rect 27448 2808 29184 2836
rect 29178 2796 29184 2808
rect 29236 2796 29242 2848
rect 30006 2796 30012 2848
rect 30064 2836 30070 2848
rect 30374 2836 30380 2848
rect 30064 2808 30380 2836
rect 30064 2796 30070 2808
rect 30374 2796 30380 2808
rect 30432 2796 30438 2848
rect 32766 2796 32772 2848
rect 32824 2836 32830 2848
rect 34054 2836 34060 2848
rect 32824 2808 34060 2836
rect 32824 2796 32830 2808
rect 34054 2796 34060 2808
rect 34112 2796 34118 2848
rect 36170 2836 36176 2848
rect 36131 2808 36176 2836
rect 36170 2796 36176 2808
rect 36228 2796 36234 2848
rect 36906 2796 36912 2848
rect 36964 2836 36970 2848
rect 39209 2839 39267 2845
rect 39209 2836 39221 2839
rect 36964 2808 39221 2836
rect 36964 2796 36970 2808
rect 39209 2805 39221 2808
rect 39255 2805 39267 2839
rect 39209 2799 39267 2805
rect 41874 2796 41880 2848
rect 41932 2836 41938 2848
rect 43257 2839 43315 2845
rect 43257 2836 43269 2839
rect 41932 2808 43269 2836
rect 41932 2796 41938 2808
rect 43257 2805 43269 2808
rect 43303 2805 43315 2839
rect 43257 2799 43315 2805
rect 43530 2796 43536 2848
rect 43588 2836 43594 2848
rect 44545 2839 44603 2845
rect 44545 2836 44557 2839
rect 43588 2808 44557 2836
rect 43588 2796 43594 2808
rect 44545 2805 44557 2808
rect 44591 2805 44603 2839
rect 44545 2799 44603 2805
rect 44910 2796 44916 2848
rect 44968 2836 44974 2848
rect 45833 2839 45891 2845
rect 45833 2836 45845 2839
rect 44968 2808 45845 2836
rect 44968 2796 44974 2808
rect 45833 2805 45845 2808
rect 45879 2805 45891 2839
rect 45833 2799 45891 2805
rect 46290 2796 46296 2848
rect 46348 2836 46354 2848
rect 47121 2839 47179 2845
rect 47121 2836 47133 2839
rect 46348 2808 47133 2836
rect 46348 2796 46354 2808
rect 47121 2805 47133 2808
rect 47167 2805 47179 2839
rect 47121 2799 47179 2805
rect 48498 2796 48504 2848
rect 48556 2836 48562 2848
rect 49237 2839 49295 2845
rect 49237 2836 49249 2839
rect 48556 2808 49249 2836
rect 48556 2796 48562 2808
rect 49237 2805 49249 2808
rect 49283 2805 49295 2839
rect 49237 2799 49295 2805
rect 49602 2796 49608 2848
rect 49660 2836 49666 2848
rect 50525 2839 50583 2845
rect 50525 2836 50537 2839
rect 49660 2808 50537 2836
rect 49660 2796 49666 2808
rect 50525 2805 50537 2808
rect 50571 2805 50583 2839
rect 50525 2799 50583 2805
rect 50614 2796 50620 2848
rect 50672 2836 50678 2848
rect 51169 2839 51227 2845
rect 51169 2836 51181 2839
rect 50672 2808 51181 2836
rect 50672 2796 50678 2808
rect 51169 2805 51181 2808
rect 51215 2805 51227 2839
rect 51169 2799 51227 2805
rect 51534 2796 51540 2848
rect 51592 2836 51598 2848
rect 52457 2839 52515 2845
rect 52457 2836 52469 2839
rect 51592 2808 52469 2836
rect 51592 2796 51598 2808
rect 52457 2805 52469 2808
rect 52503 2805 52515 2839
rect 52457 2799 52515 2805
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 22465 2635 22523 2641
rect 22465 2601 22477 2635
rect 22511 2632 22523 2635
rect 23566 2632 23572 2644
rect 22511 2604 23572 2632
rect 22511 2601 22523 2604
rect 22465 2595 22523 2601
rect 23566 2592 23572 2604
rect 23624 2592 23630 2644
rect 23753 2635 23811 2641
rect 23753 2601 23765 2635
rect 23799 2632 23811 2635
rect 25590 2632 25596 2644
rect 23799 2604 25596 2632
rect 23799 2601 23811 2604
rect 23753 2595 23811 2601
rect 25590 2592 25596 2604
rect 25648 2592 25654 2644
rect 37458 2632 37464 2644
rect 37419 2604 37464 2632
rect 37458 2592 37464 2604
rect 37516 2592 37522 2644
rect 38654 2632 38660 2644
rect 38615 2604 38660 2632
rect 38654 2592 38660 2604
rect 38712 2592 38718 2644
rect 47946 2592 47952 2644
rect 48004 2632 48010 2644
rect 49789 2635 49847 2641
rect 49789 2632 49801 2635
rect 48004 2604 49801 2632
rect 48004 2592 48010 2604
rect 49789 2601 49801 2604
rect 49835 2601 49847 2635
rect 49789 2595 49847 2601
rect 9033 2567 9091 2573
rect 9033 2533 9045 2567
rect 9079 2564 9091 2567
rect 9674 2564 9680 2576
rect 9079 2536 9680 2564
rect 9079 2533 9091 2536
rect 9033 2527 9091 2533
rect 9674 2524 9680 2536
rect 9732 2524 9738 2576
rect 10689 2567 10747 2573
rect 10689 2533 10701 2567
rect 10735 2564 10747 2567
rect 11330 2564 11336 2576
rect 10735 2536 11336 2564
rect 10735 2533 10747 2536
rect 10689 2527 10747 2533
rect 11330 2524 11336 2536
rect 11388 2524 11394 2576
rect 14277 2567 14335 2573
rect 14277 2533 14289 2567
rect 14323 2564 14335 2567
rect 14918 2564 14924 2576
rect 14323 2536 14924 2564
rect 14323 2533 14335 2536
rect 14277 2527 14335 2533
rect 14918 2524 14924 2536
rect 14976 2524 14982 2576
rect 17221 2567 17279 2573
rect 17221 2533 17233 2567
rect 17267 2564 17279 2567
rect 18414 2564 18420 2576
rect 17267 2536 18420 2564
rect 17267 2533 17279 2536
rect 17221 2527 17279 2533
rect 18414 2524 18420 2536
rect 18472 2524 18478 2576
rect 18509 2567 18567 2573
rect 18509 2533 18521 2567
rect 18555 2564 18567 2567
rect 20070 2564 20076 2576
rect 18555 2536 20076 2564
rect 18555 2533 18567 2536
rect 18509 2527 18567 2533
rect 20070 2524 20076 2536
rect 20128 2524 20134 2576
rect 20809 2567 20867 2573
rect 20809 2533 20821 2567
rect 20855 2564 20867 2567
rect 25038 2564 25044 2576
rect 20855 2536 25044 2564
rect 20855 2533 20867 2536
rect 20809 2527 20867 2533
rect 25038 2524 25044 2536
rect 25096 2524 25102 2576
rect 34974 2524 34980 2576
rect 35032 2564 35038 2576
rect 38013 2567 38071 2573
rect 38013 2564 38025 2567
rect 35032 2536 38025 2564
rect 35032 2524 35038 2536
rect 38013 2533 38025 2536
rect 38059 2533 38071 2567
rect 38013 2527 38071 2533
rect 38286 2524 38292 2576
rect 38344 2564 38350 2576
rect 40957 2567 41015 2573
rect 40957 2564 40969 2567
rect 38344 2536 40969 2564
rect 38344 2524 38350 2536
rect 40957 2533 40969 2536
rect 41003 2533 41015 2567
rect 40957 2527 41015 2533
rect 41598 2524 41604 2576
rect 41656 2564 41662 2576
rect 43257 2567 43315 2573
rect 43257 2564 43269 2567
rect 41656 2536 43269 2564
rect 41656 2524 41662 2536
rect 43257 2533 43269 2536
rect 43303 2533 43315 2567
rect 43257 2527 43315 2533
rect 45186 2524 45192 2576
rect 45244 2564 45250 2576
rect 46845 2567 46903 2573
rect 46845 2564 46857 2567
rect 45244 2536 46857 2564
rect 45244 2524 45250 2536
rect 46845 2533 46857 2536
rect 46891 2533 46903 2567
rect 46845 2527 46903 2533
rect 48774 2524 48780 2576
rect 48832 2564 48838 2576
rect 50433 2567 50491 2573
rect 50433 2564 50445 2567
rect 48832 2536 50445 2564
rect 48832 2524 48838 2536
rect 50433 2533 50445 2536
rect 50479 2533 50491 2567
rect 50433 2527 50491 2533
rect 50706 2524 50712 2576
rect 50764 2564 50770 2576
rect 52089 2567 52147 2573
rect 52089 2564 52101 2567
rect 50764 2536 52101 2564
rect 50764 2524 50770 2536
rect 52089 2533 52101 2536
rect 52135 2533 52147 2567
rect 52089 2527 52147 2533
rect 11977 2499 12035 2505
rect 11977 2465 11989 2499
rect 12023 2496 12035 2499
rect 12710 2496 12716 2508
rect 12023 2468 12716 2496
rect 12023 2465 12035 2468
rect 11977 2459 12035 2465
rect 12710 2456 12716 2468
rect 12768 2456 12774 2508
rect 16577 2499 16635 2505
rect 16577 2465 16589 2499
rect 16623 2496 16635 2499
rect 17586 2496 17592 2508
rect 16623 2468 17592 2496
rect 16623 2465 16635 2468
rect 16577 2459 16635 2465
rect 17586 2456 17592 2468
rect 17644 2456 17650 2508
rect 17865 2499 17923 2505
rect 17865 2465 17877 2499
rect 17911 2496 17923 2499
rect 19242 2496 19248 2508
rect 17911 2468 19248 2496
rect 17911 2465 17923 2468
rect 17865 2459 17923 2465
rect 19242 2456 19248 2468
rect 19300 2456 19306 2508
rect 19521 2499 19579 2505
rect 19521 2465 19533 2499
rect 19567 2496 19579 2499
rect 22830 2496 22836 2508
rect 19567 2468 22836 2496
rect 19567 2465 19579 2468
rect 19521 2459 19579 2465
rect 22830 2456 22836 2468
rect 22888 2456 22894 2508
rect 23109 2499 23167 2505
rect 23109 2465 23121 2499
rect 23155 2496 23167 2499
rect 25501 2499 25559 2505
rect 25501 2496 25513 2499
rect 23155 2468 25513 2496
rect 23155 2465 23167 2468
rect 23109 2459 23167 2465
rect 25501 2465 25513 2468
rect 25547 2465 25559 2499
rect 25501 2459 25559 2465
rect 27614 2456 27620 2508
rect 27672 2496 27678 2508
rect 28445 2499 28503 2505
rect 28445 2496 28457 2499
rect 27672 2468 28457 2496
rect 27672 2456 27678 2468
rect 28445 2465 28457 2468
rect 28491 2465 28503 2499
rect 29454 2496 29460 2508
rect 29415 2468 29460 2496
rect 28445 2459 28503 2465
rect 29454 2456 29460 2468
rect 29512 2456 29518 2508
rect 31110 2496 31116 2508
rect 31071 2468 31116 2496
rect 31110 2456 31116 2468
rect 31168 2456 31174 2508
rect 31754 2456 31760 2508
rect 31812 2496 31818 2508
rect 32493 2499 32551 2505
rect 32493 2496 32505 2499
rect 31812 2468 32505 2496
rect 31812 2456 31818 2468
rect 32493 2465 32505 2468
rect 32539 2465 32551 2499
rect 32493 2459 32551 2465
rect 32677 2499 32735 2505
rect 32677 2465 32689 2499
rect 32723 2496 32735 2499
rect 36170 2496 36176 2508
rect 32723 2468 36176 2496
rect 32723 2465 32735 2468
rect 32677 2459 32735 2465
rect 36170 2456 36176 2468
rect 36228 2456 36234 2508
rect 39114 2456 39120 2508
rect 39172 2496 39178 2508
rect 39172 2468 41644 2496
rect 39172 2456 39178 2468
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2428 7803 2431
rect 8202 2428 8208 2440
rect 7791 2400 8208 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8938 2428 8944 2440
rect 8435 2400 8944 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2428 9735 2431
rect 10226 2428 10232 2440
rect 9723 2400 10232 2428
rect 9723 2397 9735 2400
rect 9677 2391 9735 2397
rect 10226 2388 10232 2400
rect 10284 2388 10290 2440
rect 11333 2431 11391 2437
rect 11333 2397 11345 2431
rect 11379 2428 11391 2431
rect 11882 2428 11888 2440
rect 11379 2400 11888 2428
rect 11379 2397 11391 2400
rect 11333 2391 11391 2397
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2428 12679 2431
rect 13262 2428 13268 2440
rect 12667 2400 13268 2428
rect 12667 2397 12679 2400
rect 12621 2391 12679 2397
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 13633 2431 13691 2437
rect 13633 2397 13645 2431
rect 13679 2428 13691 2431
rect 14090 2428 14096 2440
rect 13679 2400 14096 2428
rect 13679 2397 13691 2400
rect 13633 2391 13691 2397
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 15565 2431 15623 2437
rect 15565 2397 15577 2431
rect 15611 2428 15623 2431
rect 16298 2428 16304 2440
rect 15611 2400 16304 2428
rect 15611 2397 15623 2400
rect 15565 2391 15623 2397
rect 14936 2360 14964 2391
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 20165 2431 20223 2437
rect 20165 2397 20177 2431
rect 20211 2397 20223 2431
rect 20165 2391 20223 2397
rect 21453 2431 21511 2437
rect 21453 2397 21465 2431
rect 21499 2428 21511 2431
rect 24118 2428 24124 2440
rect 21499 2400 24124 2428
rect 21499 2397 21511 2400
rect 21453 2391 21511 2397
rect 15746 2360 15752 2372
rect 14936 2332 15752 2360
rect 15746 2320 15752 2332
rect 15804 2320 15810 2372
rect 20180 2360 20208 2391
rect 24118 2388 24124 2400
rect 24176 2388 24182 2440
rect 24210 2388 24216 2440
rect 24268 2428 24274 2440
rect 35621 2431 35679 2437
rect 24268 2400 24313 2428
rect 24268 2388 24274 2400
rect 35621 2397 35633 2431
rect 35667 2428 35679 2431
rect 36538 2428 36544 2440
rect 35667 2400 36544 2428
rect 35667 2397 35679 2400
rect 35621 2391 35679 2397
rect 36538 2388 36544 2400
rect 36596 2388 36602 2440
rect 36722 2388 36728 2440
rect 36780 2428 36786 2440
rect 41616 2437 41644 2468
rect 42150 2456 42156 2508
rect 42208 2496 42214 2508
rect 43901 2499 43959 2505
rect 43901 2496 43913 2499
rect 42208 2468 43913 2496
rect 42208 2456 42214 2468
rect 43901 2465 43913 2468
rect 43947 2465 43959 2499
rect 43901 2459 43959 2465
rect 44634 2456 44640 2508
rect 44692 2496 44698 2508
rect 46201 2499 46259 2505
rect 46201 2496 46213 2499
rect 44692 2468 46213 2496
rect 44692 2456 44698 2468
rect 46201 2465 46213 2468
rect 46247 2465 46259 2499
rect 46201 2459 46259 2465
rect 47118 2456 47124 2508
rect 47176 2496 47182 2508
rect 48501 2499 48559 2505
rect 48501 2496 48513 2499
rect 47176 2468 48513 2496
rect 47176 2456 47182 2468
rect 48501 2465 48513 2468
rect 48547 2465 48559 2499
rect 48501 2459 48559 2465
rect 49878 2456 49884 2508
rect 49936 2496 49942 2508
rect 51445 2499 51503 2505
rect 51445 2496 51457 2499
rect 49936 2468 51457 2496
rect 49936 2456 49942 2468
rect 51445 2465 51457 2468
rect 51491 2465 51503 2499
rect 51445 2459 51503 2465
rect 51810 2456 51816 2508
rect 51868 2496 51874 2508
rect 53377 2499 53435 2505
rect 53377 2496 53389 2499
rect 51868 2468 53389 2496
rect 51868 2456 51874 2468
rect 53377 2465 53389 2468
rect 53423 2465 53435 2499
rect 53377 2459 53435 2465
rect 36909 2431 36967 2437
rect 36909 2428 36921 2431
rect 36780 2400 36921 2428
rect 36780 2388 36786 2400
rect 36909 2397 36921 2400
rect 36955 2428 36967 2431
rect 37369 2431 37427 2437
rect 37369 2428 37381 2431
rect 36955 2400 37381 2428
rect 36955 2397 36967 2400
rect 36909 2391 36967 2397
rect 37369 2397 37381 2400
rect 37415 2397 37427 2431
rect 39669 2431 39727 2437
rect 39669 2428 39681 2431
rect 37369 2391 37427 2397
rect 37476 2400 39681 2428
rect 23750 2360 23756 2372
rect 20180 2332 23756 2360
rect 23750 2320 23756 2332
rect 23808 2320 23814 2372
rect 24026 2320 24032 2372
rect 24084 2360 24090 2372
rect 25685 2363 25743 2369
rect 25685 2360 25697 2363
rect 24084 2332 25697 2360
rect 24084 2320 24090 2332
rect 25685 2329 25697 2332
rect 25731 2329 25743 2363
rect 25685 2323 25743 2329
rect 27246 2320 27252 2372
rect 27304 2360 27310 2372
rect 27341 2363 27399 2369
rect 27341 2360 27353 2363
rect 27304 2332 27353 2360
rect 27304 2320 27310 2332
rect 27341 2329 27353 2332
rect 27387 2329 27399 2363
rect 27341 2323 27399 2329
rect 28629 2363 28687 2369
rect 28629 2329 28641 2363
rect 28675 2329 28687 2363
rect 28629 2323 28687 2329
rect 24305 2295 24363 2301
rect 24305 2261 24317 2295
rect 24351 2292 24363 2295
rect 28644 2292 28672 2323
rect 33594 2320 33600 2372
rect 33652 2360 33658 2372
rect 33781 2363 33839 2369
rect 33781 2360 33793 2363
rect 33652 2332 33793 2360
rect 33652 2320 33658 2332
rect 33781 2329 33793 2332
rect 33827 2329 33839 2363
rect 33781 2323 33839 2329
rect 35437 2363 35495 2369
rect 35437 2329 35449 2363
rect 35483 2360 35495 2363
rect 36817 2363 36875 2369
rect 36817 2360 36829 2363
rect 35483 2332 36829 2360
rect 35483 2329 35495 2332
rect 35437 2323 35495 2329
rect 36817 2329 36829 2332
rect 36863 2329 36875 2363
rect 36817 2323 36875 2329
rect 24351 2264 28672 2292
rect 24351 2261 24363 2264
rect 24305 2255 24363 2261
rect 36354 2252 36360 2304
rect 36412 2292 36418 2304
rect 37476 2292 37504 2400
rect 39669 2397 39681 2400
rect 39715 2397 39727 2431
rect 39669 2391 39727 2397
rect 40313 2431 40371 2437
rect 40313 2397 40325 2431
rect 40359 2397 40371 2431
rect 40313 2391 40371 2397
rect 41601 2431 41659 2437
rect 41601 2397 41613 2431
rect 41647 2397 41659 2431
rect 41601 2391 41659 2397
rect 42613 2431 42671 2437
rect 42613 2397 42625 2431
rect 42659 2397 42671 2431
rect 42613 2391 42671 2397
rect 37734 2320 37740 2372
rect 37792 2360 37798 2372
rect 40328 2360 40356 2391
rect 37792 2332 40356 2360
rect 37792 2320 37798 2332
rect 40494 2320 40500 2372
rect 40552 2360 40558 2372
rect 42628 2360 42656 2391
rect 42702 2388 42708 2440
rect 42760 2428 42766 2440
rect 44545 2431 44603 2437
rect 44545 2428 44557 2431
rect 42760 2400 44557 2428
rect 42760 2388 42766 2400
rect 44545 2397 44557 2400
rect 44591 2397 44603 2431
rect 44545 2391 44603 2397
rect 45557 2431 45615 2437
rect 45557 2397 45569 2431
rect 45603 2397 45615 2431
rect 45557 2391 45615 2397
rect 40552 2332 42656 2360
rect 40552 2320 40558 2332
rect 43806 2320 43812 2372
rect 43864 2360 43870 2372
rect 45572 2360 45600 2391
rect 45738 2388 45744 2440
rect 45796 2428 45802 2440
rect 47489 2431 47547 2437
rect 47489 2428 47501 2431
rect 45796 2400 47501 2428
rect 45796 2388 45802 2400
rect 47489 2397 47501 2400
rect 47535 2397 47547 2431
rect 47489 2391 47547 2397
rect 49145 2431 49203 2437
rect 49145 2397 49157 2431
rect 49191 2397 49203 2431
rect 49145 2391 49203 2397
rect 52733 2431 52791 2437
rect 52733 2397 52745 2431
rect 52779 2397 52791 2431
rect 52733 2391 52791 2397
rect 43864 2332 45600 2360
rect 43864 2320 43870 2332
rect 47394 2320 47400 2372
rect 47452 2360 47458 2372
rect 49160 2360 49188 2391
rect 47452 2332 49188 2360
rect 47452 2320 47458 2332
rect 51258 2320 51264 2372
rect 51316 2360 51322 2372
rect 52748 2360 52776 2391
rect 51316 2332 52776 2360
rect 51316 2320 51322 2332
rect 36412 2264 37504 2292
rect 36412 2252 36418 2264
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 24118 2048 24124 2100
rect 24176 2088 24182 2100
rect 25866 2088 25872 2100
rect 24176 2060 25872 2088
rect 24176 2048 24182 2060
rect 25866 2048 25872 2060
rect 25924 2048 25930 2100
rect 23750 1368 23756 1420
rect 23808 1408 23814 1420
rect 24486 1408 24492 1420
rect 23808 1380 24492 1408
rect 23808 1368 23814 1380
rect 24486 1368 24492 1380
rect 24544 1368 24550 1420
<< via1 >>
rect 23204 57944 23256 57996
rect 15108 57876 15160 57928
rect 25044 57876 25096 57928
rect 12348 57808 12400 57860
rect 26976 57808 27028 57860
rect 27068 57808 27120 57860
rect 33692 57808 33744 57860
rect 23756 57740 23808 57792
rect 39948 57740 40000 57792
rect 41420 57740 41472 57792
rect 45192 57740 45244 57792
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 3700 57579 3752 57588
rect 3700 57545 3709 57579
rect 3709 57545 3743 57579
rect 3743 57545 3752 57579
rect 3700 57536 3752 57545
rect 5080 57536 5132 57588
rect 10600 57536 10652 57588
rect 11980 57536 12032 57588
rect 13360 57536 13412 57588
rect 14740 57536 14792 57588
rect 16120 57536 16172 57588
rect 17500 57536 17552 57588
rect 18880 57536 18932 57588
rect 20260 57536 20312 57588
rect 22100 57579 22152 57588
rect 22100 57545 22109 57579
rect 22109 57545 22143 57579
rect 22143 57545 22152 57579
rect 22100 57536 22152 57545
rect 23020 57536 23072 57588
rect 24860 57536 24912 57588
rect 25780 57536 25832 57588
rect 27160 57536 27212 57588
rect 28540 57536 28592 57588
rect 33140 57536 33192 57588
rect 35624 57536 35676 57588
rect 39948 57536 40000 57588
rect 5448 57443 5500 57452
rect 5448 57409 5457 57443
rect 5457 57409 5491 57443
rect 5491 57409 5500 57443
rect 5448 57400 5500 57409
rect 6000 57400 6052 57452
rect 6460 57400 6512 57452
rect 7380 57400 7432 57452
rect 7840 57400 7892 57452
rect 8760 57400 8812 57452
rect 9220 57400 9272 57452
rect 10968 57443 11020 57452
rect 10968 57409 10977 57443
rect 10977 57409 11011 57443
rect 11011 57409 11020 57443
rect 10968 57400 11020 57409
rect 11520 57400 11572 57452
rect 12348 57443 12400 57452
rect 12348 57409 12357 57443
rect 12357 57409 12391 57443
rect 12391 57409 12400 57443
rect 12348 57400 12400 57409
rect 14280 57400 14332 57452
rect 15108 57443 15160 57452
rect 15108 57409 15117 57443
rect 15117 57409 15151 57443
rect 15151 57409 15160 57443
rect 15108 57400 15160 57409
rect 16488 57443 16540 57452
rect 16488 57409 16497 57443
rect 16497 57409 16531 57443
rect 16531 57409 16540 57443
rect 16488 57400 16540 57409
rect 17040 57400 17092 57452
rect 17868 57443 17920 57452
rect 17868 57409 17877 57443
rect 17877 57409 17911 57443
rect 17911 57409 17920 57443
rect 17868 57400 17920 57409
rect 18420 57400 18472 57452
rect 5356 57264 5408 57316
rect 20628 57443 20680 57452
rect 20628 57409 20649 57443
rect 20649 57409 20680 57443
rect 20628 57400 20680 57409
rect 22284 57443 22336 57452
rect 22284 57409 22293 57443
rect 22293 57409 22327 57443
rect 22327 57409 22336 57443
rect 22284 57400 22336 57409
rect 23388 57443 23440 57452
rect 23388 57409 23397 57443
rect 23397 57409 23431 57443
rect 23431 57409 23440 57443
rect 24032 57443 24084 57452
rect 23388 57400 23440 57409
rect 24032 57409 24041 57443
rect 24041 57409 24075 57443
rect 24075 57409 24084 57443
rect 24032 57400 24084 57409
rect 24124 57400 24176 57452
rect 25596 57400 25648 57452
rect 21456 57307 21508 57316
rect 21456 57273 21465 57307
rect 21465 57273 21499 57307
rect 21499 57273 21508 57307
rect 21456 57264 21508 57273
rect 23940 57332 23992 57384
rect 23388 57264 23440 57316
rect 24308 57332 24360 57384
rect 24584 57332 24636 57384
rect 27160 57443 27212 57452
rect 27160 57409 27169 57443
rect 27169 57409 27203 57443
rect 27203 57409 27212 57443
rect 27160 57400 27212 57409
rect 27804 57400 27856 57452
rect 26332 57332 26384 57384
rect 29092 57400 29144 57452
rect 29552 57468 29604 57520
rect 42156 57536 42208 57588
rect 43352 57536 43404 57588
rect 30380 57400 30432 57452
rect 30840 57400 30892 57452
rect 31300 57332 31352 57384
rect 20628 57196 20680 57248
rect 23848 57239 23900 57248
rect 23848 57205 23857 57239
rect 23857 57205 23891 57239
rect 23891 57205 23900 57239
rect 23848 57196 23900 57205
rect 29184 57264 29236 57316
rect 31760 57400 31812 57452
rect 45560 57468 45612 57520
rect 32772 57400 32824 57452
rect 33600 57400 33652 57452
rect 32404 57375 32456 57384
rect 32404 57341 32413 57375
rect 32413 57341 32447 57375
rect 32447 57341 32456 57375
rect 32404 57332 32456 57341
rect 32956 57332 33008 57384
rect 34244 57443 34296 57452
rect 34244 57409 34253 57443
rect 34253 57409 34287 57443
rect 34287 57409 34296 57443
rect 34244 57400 34296 57409
rect 34520 57400 34572 57452
rect 34704 57400 34756 57452
rect 35624 57443 35676 57452
rect 35624 57409 35633 57443
rect 35633 57409 35667 57443
rect 35667 57409 35676 57443
rect 35624 57400 35676 57409
rect 35808 57400 35860 57452
rect 35900 57400 35952 57452
rect 37188 57400 37240 57452
rect 37280 57400 37332 57452
rect 38476 57400 38528 57452
rect 40684 57400 40736 57452
rect 25688 57196 25740 57248
rect 27160 57196 27212 57248
rect 27436 57196 27488 57248
rect 27528 57196 27580 57248
rect 28816 57196 28868 57248
rect 34336 57332 34388 57384
rect 34612 57332 34664 57384
rect 40224 57375 40276 57384
rect 33048 57196 33100 57248
rect 33324 57196 33376 57248
rect 34244 57196 34296 57248
rect 34796 57239 34848 57248
rect 34796 57205 34805 57239
rect 34805 57205 34839 57239
rect 34839 57205 34848 57239
rect 34796 57196 34848 57205
rect 35532 57196 35584 57248
rect 40224 57341 40233 57375
rect 40233 57341 40267 57375
rect 40267 57341 40276 57375
rect 40224 57332 40276 57341
rect 40500 57375 40552 57384
rect 40500 57341 40509 57375
rect 40509 57341 40543 57375
rect 40543 57341 40552 57375
rect 42800 57400 42852 57452
rect 44088 57400 44140 57452
rect 40500 57332 40552 57341
rect 43076 57332 43128 57384
rect 43352 57332 43404 57384
rect 45468 57400 45520 57452
rect 46940 57400 46992 57452
rect 48320 57400 48372 57452
rect 49700 57400 49752 57452
rect 45008 57332 45060 57384
rect 47492 57332 47544 57384
rect 43996 57264 44048 57316
rect 52460 57468 52512 57520
rect 51080 57400 51132 57452
rect 52920 57400 52972 57452
rect 53840 57400 53892 57452
rect 54208 57400 54260 57452
rect 55220 57400 55272 57452
rect 55680 57400 55732 57452
rect 40224 57196 40276 57248
rect 41052 57239 41104 57248
rect 41052 57205 41061 57239
rect 41061 57205 41095 57239
rect 41095 57205 41104 57239
rect 41052 57196 41104 57205
rect 41696 57239 41748 57248
rect 41696 57205 41705 57239
rect 41705 57205 41739 57239
rect 41739 57205 41748 57239
rect 41696 57196 41748 57205
rect 44180 57239 44232 57248
rect 44180 57205 44189 57239
rect 44189 57205 44223 57239
rect 44223 57205 44232 57239
rect 44180 57196 44232 57205
rect 44824 57239 44876 57248
rect 44824 57205 44833 57239
rect 44833 57205 44867 57239
rect 44867 57205 44876 57239
rect 44824 57196 44876 57205
rect 44916 57196 44968 57248
rect 46388 57239 46440 57248
rect 46388 57205 46397 57239
rect 46397 57205 46431 57239
rect 46431 57205 46440 57239
rect 46388 57196 46440 57205
rect 51632 57239 51684 57248
rect 51632 57205 51641 57239
rect 51641 57205 51675 57239
rect 51675 57205 51684 57239
rect 51632 57196 51684 57205
rect 52736 57239 52788 57248
rect 52736 57205 52745 57239
rect 52745 57205 52779 57239
rect 52779 57205 52788 57239
rect 52736 57196 52788 57205
rect 55404 57239 55456 57248
rect 55404 57205 55413 57239
rect 55413 57205 55447 57239
rect 55447 57205 55456 57239
rect 55404 57196 55456 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 4620 56992 4672 57044
rect 10140 56992 10192 57044
rect 12900 56992 12952 57044
rect 15660 56992 15712 57044
rect 19984 56992 20036 57044
rect 21180 56992 21232 57044
rect 10968 56924 11020 56976
rect 23204 56992 23256 57044
rect 23480 57035 23532 57044
rect 23480 57001 23489 57035
rect 23489 57001 23523 57035
rect 23523 57001 23532 57035
rect 23480 56992 23532 57001
rect 24124 56992 24176 57044
rect 24584 57035 24636 57044
rect 24584 57001 24593 57035
rect 24593 57001 24627 57035
rect 24627 57001 24636 57035
rect 24584 56992 24636 57001
rect 25044 57035 25096 57044
rect 25044 57001 25053 57035
rect 25053 57001 25087 57035
rect 25087 57001 25096 57035
rect 25044 56992 25096 57001
rect 27804 56992 27856 57044
rect 29092 57035 29144 57044
rect 29092 57001 29101 57035
rect 29101 57001 29135 57035
rect 29135 57001 29144 57035
rect 29092 56992 29144 57001
rect 29184 56992 29236 57044
rect 32680 56992 32732 57044
rect 40500 56992 40552 57044
rect 40776 56992 40828 57044
rect 25320 56924 25372 56976
rect 28172 56924 28224 56976
rect 28908 56924 28960 56976
rect 16488 56856 16540 56908
rect 26884 56856 26936 56908
rect 26976 56856 27028 56908
rect 23388 56831 23440 56840
rect 23388 56797 23397 56831
rect 23397 56797 23431 56831
rect 23431 56797 23440 56831
rect 23388 56788 23440 56797
rect 24032 56788 24084 56840
rect 25412 56788 25464 56840
rect 25596 56831 25648 56840
rect 25596 56797 25605 56831
rect 25605 56797 25639 56831
rect 25639 56797 25648 56831
rect 25596 56788 25648 56797
rect 25688 56831 25740 56840
rect 25688 56797 25697 56831
rect 25697 56797 25731 56831
rect 25731 56797 25740 56831
rect 25688 56788 25740 56797
rect 26516 56788 26568 56840
rect 26608 56831 26660 56840
rect 26608 56797 26617 56831
rect 26617 56797 26651 56831
rect 26651 56797 26660 56831
rect 26608 56788 26660 56797
rect 27068 56788 27120 56840
rect 29184 56856 29236 56908
rect 27528 56788 27580 56840
rect 27712 56831 27764 56840
rect 27712 56797 27721 56831
rect 27721 56797 27755 56831
rect 27755 56797 27764 56831
rect 27712 56788 27764 56797
rect 5448 56652 5500 56704
rect 23756 56652 23808 56704
rect 23940 56652 23992 56704
rect 25504 56652 25556 56704
rect 26424 56652 26476 56704
rect 27344 56652 27396 56704
rect 28356 56763 28408 56772
rect 28356 56729 28365 56763
rect 28365 56729 28399 56763
rect 28399 56729 28408 56763
rect 28724 56788 28776 56840
rect 28816 56788 28868 56840
rect 29276 56831 29328 56840
rect 29276 56797 29285 56831
rect 29285 56797 29319 56831
rect 29319 56797 29328 56831
rect 29276 56788 29328 56797
rect 29552 56899 29604 56908
rect 29552 56865 29561 56899
rect 29561 56865 29595 56899
rect 29595 56865 29604 56899
rect 29552 56856 29604 56865
rect 33324 56924 33376 56976
rect 40316 56924 40368 56976
rect 30656 56856 30708 56908
rect 31116 56899 31168 56908
rect 31116 56865 31125 56899
rect 31125 56865 31159 56899
rect 31159 56865 31168 56899
rect 31116 56856 31168 56865
rect 29828 56831 29880 56840
rect 29828 56797 29837 56831
rect 29837 56797 29871 56831
rect 29871 56797 29880 56831
rect 30932 56831 30984 56840
rect 29828 56788 29880 56797
rect 30932 56797 30941 56831
rect 30941 56797 30975 56831
rect 30975 56797 30984 56831
rect 30932 56788 30984 56797
rect 31208 56831 31260 56840
rect 31208 56797 31217 56831
rect 31217 56797 31251 56831
rect 31251 56797 31260 56831
rect 31208 56788 31260 56797
rect 35716 56856 35768 56908
rect 38292 56856 38344 56908
rect 32312 56831 32364 56840
rect 32312 56797 32321 56831
rect 32321 56797 32355 56831
rect 32355 56797 32364 56831
rect 32312 56788 32364 56797
rect 32772 56788 32824 56840
rect 33048 56831 33100 56840
rect 33048 56797 33057 56831
rect 33057 56797 33091 56831
rect 33091 56797 33100 56831
rect 33048 56788 33100 56797
rect 34336 56788 34388 56840
rect 34520 56788 34572 56840
rect 35072 56788 35124 56840
rect 35532 56788 35584 56840
rect 28356 56720 28408 56729
rect 28540 56695 28592 56704
rect 28540 56661 28549 56695
rect 28549 56661 28583 56695
rect 28583 56661 28592 56695
rect 28540 56652 28592 56661
rect 29184 56652 29236 56704
rect 31760 56695 31812 56704
rect 31760 56661 31769 56695
rect 31769 56661 31803 56695
rect 31803 56661 31812 56695
rect 31760 56652 31812 56661
rect 31944 56695 31996 56704
rect 31944 56661 31953 56695
rect 31953 56661 31987 56695
rect 31987 56661 31996 56695
rect 35164 56720 35216 56772
rect 31944 56652 31996 56661
rect 33692 56652 33744 56704
rect 35072 56652 35124 56704
rect 36452 56831 36504 56840
rect 36452 56797 36461 56831
rect 36461 56797 36495 56831
rect 36495 56797 36504 56831
rect 36452 56788 36504 56797
rect 36728 56831 36780 56840
rect 36728 56797 36737 56831
rect 36737 56797 36771 56831
rect 36771 56797 36780 56831
rect 36728 56788 36780 56797
rect 37924 56831 37976 56840
rect 37924 56797 37933 56831
rect 37933 56797 37967 56831
rect 37967 56797 37976 56831
rect 37924 56788 37976 56797
rect 38108 56831 38160 56840
rect 38108 56797 38117 56831
rect 38117 56797 38151 56831
rect 38151 56797 38160 56831
rect 38108 56788 38160 56797
rect 40224 56856 40276 56908
rect 38752 56831 38804 56840
rect 38752 56797 38761 56831
rect 38761 56797 38795 56831
rect 38795 56797 38804 56831
rect 41604 56856 41656 56908
rect 38752 56788 38804 56797
rect 40684 56831 40736 56840
rect 40684 56797 40693 56831
rect 40693 56797 40727 56831
rect 40727 56797 40736 56831
rect 40684 56788 40736 56797
rect 41328 56831 41380 56856
rect 41328 56804 41334 56831
rect 41334 56804 41368 56831
rect 41368 56804 41380 56831
rect 42156 56788 42208 56840
rect 47400 56992 47452 57044
rect 48780 56992 48832 57044
rect 50160 56992 50212 57044
rect 51540 56992 51592 57044
rect 53380 56992 53432 57044
rect 54300 56992 54352 57044
rect 54760 56992 54812 57044
rect 55220 56992 55272 57044
rect 56140 56992 56192 57044
rect 43812 56967 43864 56976
rect 43812 56933 43821 56967
rect 43821 56933 43855 56967
rect 43855 56933 43864 56967
rect 43812 56924 43864 56933
rect 43904 56899 43956 56908
rect 43904 56865 43913 56899
rect 43913 56865 43947 56899
rect 43947 56865 43956 56899
rect 43904 56856 43956 56865
rect 43168 56831 43220 56840
rect 36544 56720 36596 56772
rect 41512 56720 41564 56772
rect 43168 56797 43177 56831
rect 43177 56797 43211 56831
rect 43211 56797 43220 56831
rect 43168 56788 43220 56797
rect 43996 56788 44048 56840
rect 45468 56924 45520 56976
rect 46020 56924 46072 56976
rect 49240 56924 49292 56976
rect 50620 56924 50672 56976
rect 52000 56924 52052 56976
rect 47860 56856 47912 56908
rect 45192 56831 45244 56840
rect 45192 56797 45201 56831
rect 45201 56797 45235 56831
rect 45235 56797 45244 56831
rect 45192 56788 45244 56797
rect 46204 56831 46256 56840
rect 46204 56797 46213 56831
rect 46213 56797 46247 56831
rect 46247 56797 46256 56831
rect 46204 56788 46256 56797
rect 46756 56788 46808 56840
rect 36084 56695 36136 56704
rect 36084 56661 36093 56695
rect 36093 56661 36127 56695
rect 36127 56661 36136 56695
rect 36084 56652 36136 56661
rect 36176 56652 36228 56704
rect 40316 56652 40368 56704
rect 41420 56652 41472 56704
rect 42432 56652 42484 56704
rect 42616 56652 42668 56704
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 23480 56491 23532 56500
rect 23480 56457 23489 56491
rect 23489 56457 23523 56491
rect 23523 56457 23532 56491
rect 23480 56448 23532 56457
rect 26516 56448 26568 56500
rect 26884 56491 26936 56500
rect 17868 56380 17920 56432
rect 26884 56457 26893 56491
rect 26893 56457 26927 56491
rect 26927 56457 26936 56491
rect 26884 56448 26936 56457
rect 27712 56448 27764 56500
rect 28264 56448 28316 56500
rect 29828 56448 29880 56500
rect 31208 56448 31260 56500
rect 22560 56312 22612 56364
rect 23848 56312 23900 56364
rect 25504 56355 25556 56364
rect 25504 56321 25513 56355
rect 25513 56321 25547 56355
rect 25547 56321 25556 56355
rect 25504 56312 25556 56321
rect 26240 56355 26292 56364
rect 26240 56321 26249 56355
rect 26249 56321 26283 56355
rect 26283 56321 26292 56355
rect 26240 56312 26292 56321
rect 5356 56108 5408 56160
rect 24308 56244 24360 56296
rect 24768 56244 24820 56296
rect 26976 56380 27028 56432
rect 27436 56380 27488 56432
rect 26884 56312 26936 56364
rect 27344 56355 27396 56364
rect 27344 56321 27353 56355
rect 27353 56321 27387 56355
rect 27387 56321 27396 56355
rect 27344 56312 27396 56321
rect 27620 56312 27672 56364
rect 27712 56312 27764 56364
rect 28172 56355 28224 56364
rect 28172 56321 28181 56355
rect 28181 56321 28215 56355
rect 28215 56321 28224 56355
rect 28172 56312 28224 56321
rect 28448 56312 28500 56364
rect 29276 56380 29328 56432
rect 29184 56312 29236 56364
rect 30104 56380 30156 56432
rect 32956 56380 33008 56432
rect 29920 56312 29972 56364
rect 31760 56312 31812 56364
rect 32220 56312 32272 56364
rect 34796 56448 34848 56500
rect 35164 56448 35216 56500
rect 36452 56448 36504 56500
rect 35716 56423 35768 56432
rect 33324 56355 33376 56364
rect 26332 56219 26384 56228
rect 25688 56151 25740 56160
rect 25688 56117 25697 56151
rect 25697 56117 25731 56151
rect 25731 56117 25740 56151
rect 25688 56108 25740 56117
rect 26332 56185 26341 56219
rect 26341 56185 26375 56219
rect 26375 56185 26384 56219
rect 26332 56176 26384 56185
rect 31116 56244 31168 56296
rect 31576 56244 31628 56296
rect 33324 56321 33333 56355
rect 33333 56321 33367 56355
rect 33367 56321 33376 56355
rect 33324 56312 33376 56321
rect 35716 56389 35725 56423
rect 35725 56389 35759 56423
rect 35759 56389 35768 56423
rect 35716 56380 35768 56389
rect 36820 56448 36872 56500
rect 41052 56448 41104 56500
rect 43260 56448 43312 56500
rect 46388 56448 46440 56500
rect 48320 56491 48372 56500
rect 48320 56457 48329 56491
rect 48329 56457 48363 56491
rect 48363 56457 48372 56491
rect 48320 56448 48372 56457
rect 49700 56491 49752 56500
rect 49700 56457 49709 56491
rect 49709 56457 49743 56491
rect 49743 56457 49752 56491
rect 49700 56448 49752 56457
rect 51080 56448 51132 56500
rect 52460 56491 52512 56500
rect 52460 56457 52469 56491
rect 52469 56457 52503 56491
rect 52503 56457 52512 56491
rect 52460 56448 52512 56457
rect 54208 56491 54260 56500
rect 54208 56457 54217 56491
rect 54217 56457 54251 56491
rect 54251 56457 54260 56491
rect 54208 56448 54260 56457
rect 39028 56380 39080 56432
rect 33600 56355 33652 56364
rect 33600 56321 33609 56355
rect 33609 56321 33643 56355
rect 33643 56321 33652 56355
rect 33600 56312 33652 56321
rect 34612 56355 34664 56364
rect 33140 56244 33192 56296
rect 34612 56321 34621 56355
rect 34621 56321 34655 56355
rect 34655 56321 34664 56355
rect 34612 56312 34664 56321
rect 35532 56355 35584 56364
rect 35532 56321 35541 56355
rect 35541 56321 35575 56355
rect 35575 56321 35584 56355
rect 35532 56312 35584 56321
rect 36544 56312 36596 56364
rect 36728 56355 36780 56364
rect 36728 56321 36737 56355
rect 36737 56321 36771 56355
rect 36771 56321 36780 56355
rect 41696 56380 41748 56432
rect 43168 56380 43220 56432
rect 43352 56423 43404 56432
rect 43352 56389 43361 56423
rect 43361 56389 43395 56423
rect 43395 56389 43404 56423
rect 43352 56380 43404 56389
rect 43720 56380 43772 56432
rect 46204 56380 46256 56432
rect 36728 56312 36780 56321
rect 38568 56287 38620 56296
rect 38568 56253 38577 56287
rect 38577 56253 38611 56287
rect 38611 56253 38620 56287
rect 38568 56244 38620 56253
rect 38292 56176 38344 56228
rect 38936 56287 38988 56296
rect 38936 56253 38945 56287
rect 38945 56253 38979 56287
rect 38979 56253 38988 56287
rect 38936 56244 38988 56253
rect 40224 56355 40276 56364
rect 40224 56321 40233 56355
rect 40233 56321 40267 56355
rect 40267 56321 40276 56355
rect 40224 56312 40276 56321
rect 40868 56312 40920 56364
rect 41052 56355 41104 56364
rect 41052 56321 41061 56355
rect 41061 56321 41095 56355
rect 41095 56321 41104 56355
rect 41052 56312 41104 56321
rect 42156 56355 42208 56364
rect 42156 56321 42165 56355
rect 42165 56321 42199 56355
rect 42199 56321 42208 56355
rect 42156 56312 42208 56321
rect 42248 56355 42300 56364
rect 42248 56321 42257 56355
rect 42257 56321 42291 56355
rect 42291 56321 42300 56355
rect 42248 56312 42300 56321
rect 40500 56287 40552 56296
rect 40500 56253 40509 56287
rect 40509 56253 40543 56287
rect 40543 56253 40552 56287
rect 40500 56244 40552 56253
rect 40684 56244 40736 56296
rect 41144 56244 41196 56296
rect 41420 56244 41472 56296
rect 41604 56244 41656 56296
rect 42524 56355 42576 56364
rect 42524 56321 42533 56355
rect 42533 56321 42567 56355
rect 42567 56321 42576 56355
rect 42524 56312 42576 56321
rect 43076 56312 43128 56364
rect 43536 56355 43588 56364
rect 43536 56321 43545 56355
rect 43545 56321 43579 56355
rect 43579 56321 43588 56355
rect 43536 56312 43588 56321
rect 43996 56312 44048 56364
rect 45468 56312 45520 56364
rect 45652 56355 45704 56364
rect 45652 56321 45661 56355
rect 45661 56321 45695 56355
rect 45695 56321 45704 56355
rect 45652 56312 45704 56321
rect 46480 56312 46532 56364
rect 44548 56287 44600 56296
rect 44548 56253 44557 56287
rect 44557 56253 44591 56287
rect 44591 56253 44600 56287
rect 44548 56244 44600 56253
rect 45100 56244 45152 56296
rect 26608 56108 26660 56160
rect 27620 56108 27672 56160
rect 29552 56108 29604 56160
rect 30656 56151 30708 56160
rect 30656 56117 30665 56151
rect 30665 56117 30699 56151
rect 30699 56117 30708 56151
rect 30656 56108 30708 56117
rect 30932 56108 30984 56160
rect 31852 56151 31904 56160
rect 31852 56117 31861 56151
rect 31861 56117 31895 56151
rect 31895 56117 31904 56151
rect 31852 56108 31904 56117
rect 33048 56108 33100 56160
rect 33324 56108 33376 56160
rect 35716 56108 35768 56160
rect 36636 56108 36688 56160
rect 39856 56151 39908 56160
rect 39856 56117 39865 56151
rect 39865 56117 39899 56151
rect 39899 56117 39908 56151
rect 39856 56108 39908 56117
rect 40684 56108 40736 56160
rect 41420 56151 41472 56160
rect 41420 56117 41429 56151
rect 41429 56117 41463 56151
rect 41463 56117 41472 56151
rect 44640 56176 44692 56228
rect 41420 56108 41472 56117
rect 42892 56108 42944 56160
rect 45468 56151 45520 56160
rect 45468 56117 45477 56151
rect 45477 56117 45511 56151
rect 45511 56117 45520 56151
rect 45468 56108 45520 56117
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 25596 55904 25648 55956
rect 26332 55904 26384 55956
rect 30932 55904 30984 55956
rect 33784 55904 33836 55956
rect 36728 55904 36780 55956
rect 37924 55904 37976 55956
rect 38292 55904 38344 55956
rect 40868 55904 40920 55956
rect 42524 55904 42576 55956
rect 43168 55904 43220 55956
rect 44548 55904 44600 55956
rect 46756 55947 46808 55956
rect 26884 55836 26936 55888
rect 24768 55768 24820 55820
rect 23756 55700 23808 55752
rect 25412 55743 25464 55752
rect 25412 55709 25421 55743
rect 25421 55709 25455 55743
rect 25455 55709 25464 55743
rect 28264 55768 28316 55820
rect 28448 55811 28500 55820
rect 28448 55777 28457 55811
rect 28457 55777 28491 55811
rect 28491 55777 28500 55811
rect 28448 55768 28500 55777
rect 28540 55768 28592 55820
rect 29368 55768 29420 55820
rect 25412 55700 25464 55709
rect 24032 55607 24084 55616
rect 24032 55573 24041 55607
rect 24041 55573 24075 55607
rect 24075 55573 24084 55607
rect 24032 55564 24084 55573
rect 26976 55743 27028 55752
rect 26976 55709 26985 55743
rect 26985 55709 27019 55743
rect 27019 55709 27028 55743
rect 26976 55700 27028 55709
rect 28632 55743 28684 55752
rect 28632 55709 28641 55743
rect 28641 55709 28675 55743
rect 28675 55709 28684 55743
rect 28632 55700 28684 55709
rect 28816 55743 28868 55752
rect 28816 55709 28825 55743
rect 28825 55709 28859 55743
rect 28859 55709 28868 55743
rect 28816 55700 28868 55709
rect 29920 55768 29972 55820
rect 35532 55836 35584 55888
rect 34980 55811 35032 55820
rect 34980 55777 34989 55811
rect 34989 55777 35023 55811
rect 35023 55777 35032 55811
rect 34980 55768 35032 55777
rect 36636 55811 36688 55820
rect 36636 55777 36645 55811
rect 36645 55777 36679 55811
rect 36679 55777 36688 55811
rect 36636 55768 36688 55777
rect 38384 55836 38436 55888
rect 29736 55700 29788 55752
rect 30104 55700 30156 55752
rect 30840 55743 30892 55752
rect 30840 55709 30849 55743
rect 30849 55709 30883 55743
rect 30883 55709 30892 55743
rect 30840 55700 30892 55709
rect 31300 55743 31352 55752
rect 31300 55709 31309 55743
rect 31309 55709 31343 55743
rect 31343 55709 31352 55743
rect 31300 55700 31352 55709
rect 32404 55743 32456 55752
rect 27896 55632 27948 55684
rect 29000 55632 29052 55684
rect 30748 55632 30800 55684
rect 31116 55675 31168 55684
rect 31116 55641 31125 55675
rect 31125 55641 31159 55675
rect 31159 55641 31168 55675
rect 31116 55632 31168 55641
rect 32404 55709 32413 55743
rect 32413 55709 32447 55743
rect 32447 55709 32456 55743
rect 32404 55700 32456 55709
rect 32680 55700 32732 55752
rect 33048 55743 33100 55752
rect 33048 55709 33057 55743
rect 33057 55709 33091 55743
rect 33091 55709 33100 55743
rect 33048 55700 33100 55709
rect 33232 55743 33284 55752
rect 33232 55709 33241 55743
rect 33241 55709 33275 55743
rect 33275 55709 33284 55743
rect 33232 55700 33284 55709
rect 33692 55700 33744 55752
rect 34060 55700 34112 55752
rect 34796 55700 34848 55752
rect 32864 55675 32916 55684
rect 29276 55564 29328 55616
rect 29460 55607 29512 55616
rect 29460 55573 29469 55607
rect 29469 55573 29503 55607
rect 29503 55573 29512 55607
rect 29460 55564 29512 55573
rect 30656 55564 30708 55616
rect 32312 55607 32364 55616
rect 32312 55573 32321 55607
rect 32321 55573 32355 55607
rect 32355 55573 32364 55607
rect 32312 55564 32364 55573
rect 32864 55641 32873 55675
rect 32873 55641 32907 55675
rect 32907 55641 32916 55675
rect 32864 55632 32916 55641
rect 34336 55632 34388 55684
rect 36084 55700 36136 55752
rect 36544 55743 36596 55752
rect 36544 55709 36553 55743
rect 36553 55709 36587 55743
rect 36587 55709 36596 55743
rect 36544 55700 36596 55709
rect 37924 55700 37976 55752
rect 38292 55743 38344 55752
rect 38292 55709 38301 55743
rect 38301 55709 38335 55743
rect 38335 55709 38344 55743
rect 38292 55700 38344 55709
rect 38568 55836 38620 55888
rect 38936 55836 38988 55888
rect 40408 55836 40460 55888
rect 40776 55836 40828 55888
rect 40960 55836 41012 55888
rect 41696 55836 41748 55888
rect 42248 55836 42300 55888
rect 42800 55836 42852 55888
rect 40592 55768 40644 55820
rect 38660 55743 38712 55752
rect 38660 55709 38669 55743
rect 38669 55709 38703 55743
rect 38703 55709 38712 55743
rect 39304 55743 39356 55752
rect 38660 55700 38712 55709
rect 39304 55709 39313 55743
rect 39313 55709 39347 55743
rect 39347 55709 39356 55743
rect 39304 55700 39356 55709
rect 39488 55743 39540 55752
rect 39488 55709 39497 55743
rect 39497 55709 39531 55743
rect 39531 55709 39540 55743
rect 39488 55700 39540 55709
rect 39948 55700 40000 55752
rect 39120 55675 39172 55684
rect 35164 55564 35216 55616
rect 39120 55641 39129 55675
rect 39129 55641 39163 55675
rect 39163 55641 39172 55675
rect 39120 55632 39172 55641
rect 40408 55675 40460 55684
rect 40408 55641 40417 55675
rect 40417 55641 40451 55675
rect 40451 55641 40460 55675
rect 40408 55632 40460 55641
rect 40592 55675 40644 55684
rect 40592 55641 40601 55675
rect 40601 55641 40635 55675
rect 40635 55641 40644 55675
rect 40592 55632 40644 55641
rect 40868 55700 40920 55752
rect 42616 55700 42668 55752
rect 42800 55743 42852 55752
rect 42800 55709 42809 55743
rect 42809 55709 42843 55743
rect 42843 55709 42852 55743
rect 42800 55700 42852 55709
rect 41328 55632 41380 55684
rect 44272 55836 44324 55888
rect 46756 55913 46765 55947
rect 46765 55913 46799 55947
rect 46799 55913 46808 55947
rect 46756 55904 46808 55913
rect 46940 55904 46992 55956
rect 45008 55879 45060 55888
rect 45008 55845 45017 55879
rect 45017 55845 45051 55879
rect 45051 55845 45060 55879
rect 45008 55836 45060 55845
rect 45652 55836 45704 55888
rect 55404 55836 55456 55888
rect 43536 55768 43588 55820
rect 43996 55743 44048 55752
rect 43996 55709 44005 55743
rect 44005 55709 44039 55743
rect 44039 55709 44048 55743
rect 43996 55700 44048 55709
rect 44548 55700 44600 55752
rect 47492 55768 47544 55820
rect 44916 55743 44968 55752
rect 44916 55709 44925 55743
rect 44925 55709 44959 55743
rect 44959 55709 44968 55743
rect 44916 55700 44968 55709
rect 44732 55632 44784 55684
rect 45468 55700 45520 55752
rect 38108 55564 38160 55616
rect 40684 55564 40736 55616
rect 40776 55564 40828 55616
rect 42892 55564 42944 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 23388 55360 23440 55412
rect 25780 55360 25832 55412
rect 26240 55403 26292 55412
rect 26240 55369 26249 55403
rect 26249 55369 26283 55403
rect 26283 55369 26292 55403
rect 26240 55360 26292 55369
rect 28356 55360 28408 55412
rect 28816 55360 28868 55412
rect 30748 55403 30800 55412
rect 29460 55292 29512 55344
rect 24032 55267 24084 55276
rect 24032 55233 24041 55267
rect 24041 55233 24075 55267
rect 24075 55233 24084 55267
rect 24032 55224 24084 55233
rect 25688 55267 25740 55276
rect 25688 55233 25697 55267
rect 25697 55233 25731 55267
rect 25731 55233 25740 55267
rect 25688 55224 25740 55233
rect 26424 55267 26476 55276
rect 26424 55233 26433 55267
rect 26433 55233 26467 55267
rect 26467 55233 26476 55267
rect 26424 55224 26476 55233
rect 26608 55224 26660 55276
rect 27528 55267 27580 55276
rect 27528 55233 27537 55267
rect 27537 55233 27571 55267
rect 27571 55233 27580 55267
rect 27528 55224 27580 55233
rect 27712 55267 27764 55276
rect 27712 55233 27721 55267
rect 27721 55233 27755 55267
rect 27755 55233 27764 55267
rect 27712 55224 27764 55233
rect 28448 55224 28500 55276
rect 28540 55156 28592 55208
rect 30748 55369 30757 55403
rect 30757 55369 30791 55403
rect 30791 55369 30800 55403
rect 30748 55360 30800 55369
rect 31300 55360 31352 55412
rect 29736 55335 29788 55344
rect 29736 55301 29745 55335
rect 29745 55301 29779 55335
rect 29779 55301 29788 55335
rect 29920 55335 29972 55344
rect 29736 55292 29788 55301
rect 29920 55301 29929 55335
rect 29929 55301 29963 55335
rect 29963 55301 29972 55335
rect 29920 55292 29972 55301
rect 34980 55403 35032 55412
rect 33600 55335 33652 55344
rect 33600 55301 33609 55335
rect 33609 55301 33643 55335
rect 33643 55301 33652 55335
rect 33600 55292 33652 55301
rect 34336 55335 34388 55344
rect 34336 55301 34345 55335
rect 34345 55301 34379 55335
rect 34379 55301 34388 55335
rect 34336 55292 34388 55301
rect 34980 55369 34989 55403
rect 34989 55369 35023 55403
rect 35023 55369 35032 55403
rect 34980 55360 35032 55369
rect 35164 55360 35216 55412
rect 35440 55360 35492 55412
rect 36544 55360 36596 55412
rect 38384 55360 38436 55412
rect 39120 55360 39172 55412
rect 40500 55360 40552 55412
rect 40684 55360 40736 55412
rect 41236 55360 41288 55412
rect 42432 55360 42484 55412
rect 34612 55292 34664 55344
rect 30380 55267 30432 55276
rect 30380 55233 30389 55267
rect 30389 55233 30423 55267
rect 30423 55233 30432 55267
rect 30380 55224 30432 55233
rect 30564 55267 30616 55276
rect 30564 55233 30573 55267
rect 30573 55233 30607 55267
rect 30607 55233 30616 55267
rect 30564 55224 30616 55233
rect 31576 55224 31628 55276
rect 32680 55267 32732 55276
rect 32680 55233 32689 55267
rect 32689 55233 32723 55267
rect 32723 55233 32732 55267
rect 32680 55224 32732 55233
rect 32312 55156 32364 55208
rect 33324 55224 33376 55276
rect 33692 55267 33744 55276
rect 33692 55233 33701 55267
rect 33701 55233 33735 55267
rect 33735 55233 33744 55267
rect 33692 55224 33744 55233
rect 35164 55267 35216 55276
rect 35164 55233 35173 55267
rect 35173 55233 35207 55267
rect 35207 55233 35216 55267
rect 35164 55224 35216 55233
rect 35624 55292 35676 55344
rect 34428 55156 34480 55208
rect 35532 55224 35584 55276
rect 35716 55224 35768 55276
rect 34888 55088 34940 55140
rect 35716 55088 35768 55140
rect 36452 55224 36504 55276
rect 38660 55292 38712 55344
rect 39948 55335 40000 55344
rect 38384 55224 38436 55276
rect 39488 55224 39540 55276
rect 39948 55301 39957 55335
rect 39957 55301 39991 55335
rect 39991 55301 40000 55335
rect 39948 55292 40000 55301
rect 40224 55292 40276 55344
rect 44088 55360 44140 55412
rect 45192 55360 45244 55412
rect 45560 55403 45612 55412
rect 45560 55369 45569 55403
rect 45569 55369 45603 55403
rect 45603 55369 45612 55403
rect 45560 55360 45612 55369
rect 45652 55292 45704 55344
rect 39856 55267 39908 55276
rect 39856 55233 39865 55267
rect 39865 55233 39899 55267
rect 39899 55233 39908 55267
rect 39856 55224 39908 55233
rect 39304 55156 39356 55208
rect 41972 55224 42024 55276
rect 42340 55224 42392 55276
rect 41144 55156 41196 55208
rect 41880 55156 41932 55208
rect 42708 55088 42760 55140
rect 24768 55063 24820 55072
rect 24768 55029 24777 55063
rect 24777 55029 24811 55063
rect 24811 55029 24820 55063
rect 24768 55020 24820 55029
rect 27620 55063 27672 55072
rect 27620 55029 27629 55063
rect 27629 55029 27663 55063
rect 27663 55029 27672 55063
rect 27620 55020 27672 55029
rect 28448 55020 28500 55072
rect 31852 55063 31904 55072
rect 31852 55029 31861 55063
rect 31861 55029 31895 55063
rect 31895 55029 31904 55063
rect 31852 55020 31904 55029
rect 32404 55020 32456 55072
rect 37280 55020 37332 55072
rect 40316 55020 40368 55072
rect 41236 55020 41288 55072
rect 41604 55063 41656 55072
rect 41604 55029 41613 55063
rect 41613 55029 41647 55063
rect 41647 55029 41656 55063
rect 41604 55020 41656 55029
rect 41880 55063 41932 55072
rect 41880 55029 41889 55063
rect 41889 55029 41923 55063
rect 41923 55029 41932 55063
rect 41880 55020 41932 55029
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 26608 54816 26660 54868
rect 26700 54816 26752 54868
rect 28080 54816 28132 54868
rect 28724 54816 28776 54868
rect 29552 54816 29604 54868
rect 30840 54816 30892 54868
rect 34796 54816 34848 54868
rect 35348 54816 35400 54868
rect 36360 54816 36412 54868
rect 37280 54816 37332 54868
rect 37740 54816 37792 54868
rect 38476 54859 38528 54868
rect 38476 54825 38485 54859
rect 38485 54825 38519 54859
rect 38519 54825 38528 54859
rect 38476 54816 38528 54825
rect 39948 54816 40000 54868
rect 41696 54859 41748 54868
rect 41696 54825 41705 54859
rect 41705 54825 41739 54859
rect 41739 54825 41748 54859
rect 41696 54816 41748 54825
rect 45008 54816 45060 54868
rect 24768 54748 24820 54800
rect 26976 54748 27028 54800
rect 28540 54748 28592 54800
rect 30380 54748 30432 54800
rect 33876 54680 33928 54732
rect 29184 54544 29236 54596
rect 29000 54476 29052 54528
rect 29644 54655 29696 54664
rect 29644 54621 29653 54655
rect 29653 54621 29687 54655
rect 29687 54621 29696 54655
rect 29644 54612 29696 54621
rect 30380 54612 30432 54664
rect 32404 54655 32456 54664
rect 30564 54544 30616 54596
rect 31116 54544 31168 54596
rect 32404 54621 32413 54655
rect 32413 54621 32447 54655
rect 32447 54621 32456 54655
rect 32404 54612 32456 54621
rect 33140 54612 33192 54664
rect 33324 54655 33376 54664
rect 33324 54621 33333 54655
rect 33333 54621 33367 54655
rect 33367 54621 33376 54655
rect 33324 54612 33376 54621
rect 34428 54655 34480 54664
rect 34428 54621 34437 54655
rect 34437 54621 34471 54655
rect 34471 54621 34480 54655
rect 34428 54612 34480 54621
rect 35716 54680 35768 54732
rect 39488 54748 39540 54800
rect 39856 54680 39908 54732
rect 40868 54680 40920 54732
rect 34612 54655 34664 54664
rect 34612 54621 34621 54655
rect 34621 54621 34655 54655
rect 34655 54621 34664 54655
rect 39212 54655 39264 54664
rect 34612 54612 34664 54621
rect 39212 54621 39221 54655
rect 39221 54621 39255 54655
rect 39255 54621 39264 54655
rect 39212 54612 39264 54621
rect 41880 54680 41932 54732
rect 44916 54680 44968 54732
rect 41236 54655 41288 54664
rect 41236 54621 41245 54655
rect 41245 54621 41279 54655
rect 41279 54621 41288 54655
rect 41236 54612 41288 54621
rect 32588 54544 32640 54596
rect 38752 54544 38804 54596
rect 41972 54544 42024 54596
rect 42708 54655 42760 54664
rect 42708 54621 42717 54655
rect 42717 54621 42751 54655
rect 42751 54621 42760 54655
rect 42708 54612 42760 54621
rect 43536 54612 43588 54664
rect 44732 54655 44784 54664
rect 44732 54621 44741 54655
rect 44741 54621 44775 54655
rect 44775 54621 44784 54655
rect 44732 54612 44784 54621
rect 29460 54476 29512 54528
rect 32864 54519 32916 54528
rect 32864 54485 32873 54519
rect 32873 54485 32907 54519
rect 32907 54485 32916 54519
rect 32864 54476 32916 54485
rect 33508 54476 33560 54528
rect 42432 54519 42484 54528
rect 42432 54485 42441 54519
rect 42441 54485 42475 54519
rect 42475 54485 42484 54519
rect 42432 54476 42484 54485
rect 42800 54476 42852 54528
rect 44180 54476 44232 54528
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 27068 54272 27120 54324
rect 27896 54315 27948 54324
rect 27896 54281 27905 54315
rect 27905 54281 27939 54315
rect 27939 54281 27948 54315
rect 27896 54272 27948 54281
rect 28908 54315 28960 54324
rect 28908 54281 28917 54315
rect 28917 54281 28951 54315
rect 28951 54281 28960 54315
rect 28908 54272 28960 54281
rect 29184 54272 29236 54324
rect 29644 54272 29696 54324
rect 33232 54272 33284 54324
rect 33324 54272 33376 54324
rect 34612 54272 34664 54324
rect 34980 54272 35032 54324
rect 35440 54272 35492 54324
rect 36452 54272 36504 54324
rect 37188 54272 37240 54324
rect 39028 54315 39080 54324
rect 39028 54281 39037 54315
rect 39037 54281 39071 54315
rect 39071 54281 39080 54315
rect 39028 54272 39080 54281
rect 40316 54315 40368 54324
rect 40316 54281 40325 54315
rect 40325 54281 40359 54315
rect 40359 54281 40368 54315
rect 40316 54272 40368 54281
rect 41420 54272 41472 54324
rect 41972 54315 42024 54324
rect 41972 54281 41981 54315
rect 41981 54281 42015 54315
rect 42015 54281 42024 54315
rect 41972 54272 42024 54281
rect 29736 54204 29788 54256
rect 28540 54179 28592 54188
rect 28540 54145 28549 54179
rect 28549 54145 28583 54179
rect 28583 54145 28592 54179
rect 28540 54136 28592 54145
rect 32680 54204 32732 54256
rect 28448 54111 28500 54120
rect 28448 54077 28457 54111
rect 28457 54077 28491 54111
rect 28491 54077 28500 54111
rect 28448 54068 28500 54077
rect 29736 54111 29788 54120
rect 29736 54077 29745 54111
rect 29745 54077 29779 54111
rect 29779 54077 29788 54111
rect 29736 54068 29788 54077
rect 32404 54179 32456 54188
rect 32404 54145 32413 54179
rect 32413 54145 32447 54179
rect 32447 54145 32456 54179
rect 32404 54136 32456 54145
rect 34428 54136 34480 54188
rect 34980 54179 35032 54188
rect 34980 54145 35003 54179
rect 35003 54145 35032 54179
rect 35716 54179 35768 54188
rect 34980 54136 35032 54145
rect 35716 54145 35725 54179
rect 35725 54145 35759 54179
rect 35759 54145 35768 54179
rect 35716 54136 35768 54145
rect 38200 54136 38252 54188
rect 40224 54204 40276 54256
rect 42064 54204 42116 54256
rect 40040 54136 40092 54188
rect 41604 54136 41656 54188
rect 42432 54179 42484 54188
rect 26976 54000 27028 54052
rect 28632 54000 28684 54052
rect 30196 54000 30248 54052
rect 30564 54068 30616 54120
rect 32312 54111 32364 54120
rect 32312 54077 32321 54111
rect 32321 54077 32355 54111
rect 32355 54077 32364 54111
rect 32312 54068 32364 54077
rect 33876 54111 33928 54120
rect 33876 54077 33885 54111
rect 33885 54077 33919 54111
rect 33919 54077 33928 54111
rect 33876 54068 33928 54077
rect 41236 54111 41288 54120
rect 41236 54077 41245 54111
rect 41245 54077 41279 54111
rect 41279 54077 41288 54111
rect 41236 54068 41288 54077
rect 42432 54145 42441 54179
rect 42441 54145 42475 54179
rect 42475 54145 42484 54179
rect 42432 54136 42484 54145
rect 44732 54204 44784 54256
rect 42248 54068 42300 54120
rect 42616 54068 42668 54120
rect 42708 54068 42760 54120
rect 44180 54136 44232 54188
rect 45008 54136 45060 54188
rect 44916 54068 44968 54120
rect 31116 53932 31168 53984
rect 33692 53932 33744 53984
rect 34612 53932 34664 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 29000 53728 29052 53780
rect 32404 53771 32456 53780
rect 32404 53737 32413 53771
rect 32413 53737 32447 53771
rect 32447 53737 32456 53771
rect 32404 53728 32456 53737
rect 32588 53771 32640 53780
rect 32588 53737 32597 53771
rect 32597 53737 32631 53771
rect 32631 53737 32640 53771
rect 32588 53728 32640 53737
rect 33508 53771 33560 53780
rect 33508 53737 33517 53771
rect 33517 53737 33551 53771
rect 33551 53737 33560 53771
rect 33508 53728 33560 53737
rect 34888 53771 34940 53780
rect 34888 53737 34897 53771
rect 34897 53737 34931 53771
rect 34931 53737 34940 53771
rect 34888 53728 34940 53737
rect 35532 53728 35584 53780
rect 35900 53771 35952 53780
rect 35900 53737 35909 53771
rect 35909 53737 35943 53771
rect 35943 53737 35952 53771
rect 35900 53728 35952 53737
rect 40040 53728 40092 53780
rect 41880 53771 41932 53780
rect 41880 53737 41889 53771
rect 41889 53737 41923 53771
rect 41923 53737 41932 53771
rect 41880 53728 41932 53737
rect 42064 53771 42116 53780
rect 42064 53737 42073 53771
rect 42073 53737 42107 53771
rect 42107 53737 42116 53771
rect 42064 53728 42116 53737
rect 31116 53660 31168 53712
rect 33692 53660 33744 53712
rect 36452 53660 36504 53712
rect 33140 53592 33192 53644
rect 29736 53524 29788 53576
rect 30196 53567 30248 53576
rect 30196 53533 30205 53567
rect 30205 53533 30239 53567
rect 30239 53533 30248 53567
rect 30196 53524 30248 53533
rect 32864 53567 32916 53576
rect 32864 53533 32873 53567
rect 32873 53533 32907 53567
rect 32907 53533 32916 53567
rect 32864 53524 32916 53533
rect 33324 53524 33376 53576
rect 40224 53592 40276 53644
rect 40776 53635 40828 53644
rect 40776 53601 40785 53635
rect 40785 53601 40819 53635
rect 40819 53601 40828 53635
rect 40776 53592 40828 53601
rect 42248 53499 42300 53508
rect 42248 53465 42257 53499
rect 42257 53465 42291 53499
rect 42291 53465 42300 53499
rect 42248 53456 42300 53465
rect 28632 53431 28684 53440
rect 28632 53397 28641 53431
rect 28641 53397 28675 53431
rect 28675 53397 28684 53431
rect 28632 53388 28684 53397
rect 29000 53388 29052 53440
rect 42432 53388 42484 53440
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 33692 53227 33744 53236
rect 33692 53193 33701 53227
rect 33701 53193 33735 53227
rect 33735 53193 33744 53227
rect 33692 53184 33744 53193
rect 34704 53184 34756 53236
rect 40776 53227 40828 53236
rect 40776 53193 40785 53227
rect 40785 53193 40819 53227
rect 40819 53193 40828 53227
rect 40776 53184 40828 53193
rect 34888 53159 34940 53168
rect 34888 53125 34897 53159
rect 34897 53125 34931 53159
rect 34931 53125 34940 53159
rect 34888 53116 34940 53125
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 27528 52368 27580 52420
rect 34520 52368 34572 52420
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 34520 52028 34572 52080
rect 34060 51935 34112 51944
rect 34060 51901 34069 51935
rect 34069 51901 34103 51935
rect 34103 51901 34112 51935
rect 34060 51892 34112 51901
rect 35808 51935 35860 51944
rect 35808 51901 35817 51935
rect 35817 51901 35851 51935
rect 35851 51901 35860 51935
rect 35808 51892 35860 51901
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 34060 51552 34112 51604
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 29552 8440 29604 8492
rect 30196 8304 30248 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 29000 8075 29052 8084
rect 29000 8041 29009 8075
rect 29009 8041 29043 8075
rect 29043 8041 29052 8075
rect 29000 8032 29052 8041
rect 29552 7896 29604 7948
rect 29460 7871 29512 7880
rect 29460 7837 29469 7871
rect 29469 7837 29503 7871
rect 29503 7837 29512 7871
rect 29460 7828 29512 7837
rect 30012 7828 30064 7880
rect 31208 7692 31260 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 26976 7395 27028 7404
rect 26976 7361 26985 7395
rect 26985 7361 27019 7395
rect 27019 7361 27028 7395
rect 26976 7352 27028 7361
rect 29092 7352 29144 7404
rect 31576 7352 31628 7404
rect 27712 7327 27764 7336
rect 27712 7293 27721 7327
rect 27721 7293 27755 7327
rect 27755 7293 27764 7327
rect 27712 7284 27764 7293
rect 27896 7327 27948 7336
rect 27896 7293 27905 7327
rect 27905 7293 27939 7327
rect 27939 7293 27948 7327
rect 27896 7284 27948 7293
rect 29184 7327 29236 7336
rect 29184 7293 29193 7327
rect 29193 7293 29227 7327
rect 29227 7293 29236 7327
rect 29184 7284 29236 7293
rect 29552 7284 29604 7336
rect 26884 7191 26936 7200
rect 26884 7157 26893 7191
rect 26893 7157 26927 7191
rect 26927 7157 26936 7191
rect 26884 7148 26936 7157
rect 31300 7191 31352 7200
rect 31300 7157 31309 7191
rect 31309 7157 31343 7191
rect 31343 7157 31352 7191
rect 31300 7148 31352 7157
rect 33784 7148 33836 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 30564 6944 30616 6996
rect 31576 6944 31628 6996
rect 29460 6808 29512 6860
rect 30288 6851 30340 6860
rect 30288 6817 30297 6851
rect 30297 6817 30331 6851
rect 30331 6817 30340 6851
rect 30288 6808 30340 6817
rect 31208 6851 31260 6860
rect 31208 6817 31217 6851
rect 31217 6817 31251 6851
rect 31251 6817 31260 6851
rect 31208 6808 31260 6817
rect 31484 6851 31536 6860
rect 31484 6817 31493 6851
rect 31493 6817 31527 6851
rect 31527 6817 31536 6851
rect 31484 6808 31536 6817
rect 31576 6808 31628 6860
rect 26976 6740 27028 6792
rect 27620 6740 27672 6792
rect 29460 6672 29512 6724
rect 31300 6672 31352 6724
rect 26424 6647 26476 6656
rect 26424 6613 26433 6647
rect 26433 6613 26467 6647
rect 26467 6613 26476 6647
rect 26424 6604 26476 6613
rect 27804 6604 27856 6656
rect 34428 6604 34480 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 26424 6264 26476 6316
rect 29092 6400 29144 6452
rect 27804 6375 27856 6384
rect 27804 6341 27813 6375
rect 27813 6341 27847 6375
rect 27847 6341 27856 6375
rect 27804 6332 27856 6341
rect 30564 6375 30616 6384
rect 30564 6341 30573 6375
rect 30573 6341 30607 6375
rect 30607 6341 30616 6375
rect 30564 6332 30616 6341
rect 27620 6307 27672 6316
rect 27620 6273 27629 6307
rect 27629 6273 27663 6307
rect 27663 6273 27672 6307
rect 27620 6264 27672 6273
rect 29092 6264 29144 6316
rect 26976 6239 27028 6248
rect 26976 6205 26985 6239
rect 26985 6205 27019 6239
rect 27019 6205 27028 6239
rect 26976 6196 27028 6205
rect 27436 6196 27488 6248
rect 28080 6239 28132 6248
rect 28080 6205 28089 6239
rect 28089 6205 28123 6239
rect 28123 6205 28132 6239
rect 28080 6196 28132 6205
rect 32588 6239 32640 6248
rect 32588 6205 32597 6239
rect 32597 6205 32631 6239
rect 32631 6205 32640 6239
rect 32588 6196 32640 6205
rect 33048 6196 33100 6248
rect 27712 6128 27764 6180
rect 32496 6128 32548 6180
rect 25320 6103 25372 6112
rect 25320 6069 25329 6103
rect 25329 6069 25363 6103
rect 25363 6069 25372 6103
rect 25320 6060 25372 6069
rect 34244 6060 34296 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 29460 5899 29512 5908
rect 29460 5865 29469 5899
rect 29469 5865 29503 5899
rect 29503 5865 29512 5899
rect 29460 5856 29512 5865
rect 32496 5899 32548 5908
rect 32496 5865 32505 5899
rect 32505 5865 32539 5899
rect 32539 5865 32548 5899
rect 32496 5856 32548 5865
rect 33048 5899 33100 5908
rect 33048 5865 33057 5899
rect 33057 5865 33091 5899
rect 33091 5865 33100 5899
rect 33048 5856 33100 5865
rect 26424 5788 26476 5840
rect 33876 5788 33928 5840
rect 26884 5720 26936 5772
rect 27528 5763 27580 5772
rect 27528 5729 27537 5763
rect 27537 5729 27571 5763
rect 27571 5729 27580 5763
rect 27528 5720 27580 5729
rect 30012 5763 30064 5772
rect 30012 5729 30021 5763
rect 30021 5729 30055 5763
rect 30055 5729 30064 5763
rect 30012 5720 30064 5729
rect 30196 5763 30248 5772
rect 30196 5729 30205 5763
rect 30205 5729 30239 5763
rect 30239 5729 30248 5763
rect 30196 5720 30248 5729
rect 30564 5763 30616 5772
rect 30564 5729 30573 5763
rect 30573 5729 30607 5763
rect 30607 5729 30616 5763
rect 30564 5720 30616 5729
rect 30656 5720 30708 5772
rect 34244 5763 34296 5772
rect 28908 5695 28960 5704
rect 28908 5661 28917 5695
rect 28917 5661 28951 5695
rect 28951 5661 28960 5695
rect 28908 5652 28960 5661
rect 29000 5652 29052 5704
rect 29552 5695 29604 5704
rect 29552 5661 29561 5695
rect 29561 5661 29595 5695
rect 29595 5661 29604 5695
rect 29552 5652 29604 5661
rect 34244 5729 34253 5763
rect 34253 5729 34287 5763
rect 34287 5729 34296 5763
rect 34244 5720 34296 5729
rect 34428 5763 34480 5772
rect 34428 5729 34437 5763
rect 34437 5729 34471 5763
rect 34471 5729 34480 5763
rect 34428 5720 34480 5729
rect 25504 5516 25556 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 27896 5312 27948 5364
rect 25504 5287 25556 5296
rect 25504 5253 25513 5287
rect 25513 5253 25547 5287
rect 25547 5253 25556 5287
rect 25504 5244 25556 5253
rect 30840 5244 30892 5296
rect 33784 5287 33836 5296
rect 33784 5253 33793 5287
rect 33793 5253 33827 5287
rect 33827 5253 33836 5287
rect 33784 5244 33836 5253
rect 25320 5219 25372 5228
rect 25320 5185 25329 5219
rect 25329 5185 25363 5219
rect 25363 5185 25372 5219
rect 25320 5176 25372 5185
rect 27436 5176 27488 5228
rect 28908 5219 28960 5228
rect 24768 5108 24820 5160
rect 26240 5151 26292 5160
rect 26240 5117 26249 5151
rect 26249 5117 26283 5151
rect 26283 5117 26292 5151
rect 26240 5108 26292 5117
rect 26332 5040 26384 5092
rect 28908 5185 28917 5219
rect 28917 5185 28951 5219
rect 28951 5185 28960 5219
rect 28908 5176 28960 5185
rect 30380 5151 30432 5160
rect 30380 5117 30389 5151
rect 30389 5117 30423 5151
rect 30423 5117 30432 5151
rect 30380 5108 30432 5117
rect 31300 5151 31352 5160
rect 31300 5117 31309 5151
rect 31309 5117 31343 5151
rect 31343 5117 31352 5151
rect 31300 5108 31352 5117
rect 31760 5151 31812 5160
rect 31760 5117 31769 5151
rect 31769 5117 31803 5151
rect 31803 5117 31812 5151
rect 31760 5108 31812 5117
rect 33600 5151 33652 5160
rect 33600 5117 33609 5151
rect 33609 5117 33643 5151
rect 33643 5117 33652 5151
rect 33600 5108 33652 5117
rect 34060 5151 34112 5160
rect 34060 5117 34069 5151
rect 34069 5117 34103 5151
rect 34103 5117 34112 5151
rect 34060 5108 34112 5117
rect 29000 5040 29052 5092
rect 23112 4972 23164 5024
rect 25872 4972 25924 5024
rect 36084 5015 36136 5024
rect 36084 4981 36093 5015
rect 36093 4981 36127 5015
rect 36127 4981 36136 5015
rect 36084 4972 36136 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 27896 4768 27948 4820
rect 33600 4768 33652 4820
rect 23940 4700 23992 4752
rect 27252 4700 27304 4752
rect 25872 4675 25924 4684
rect 25872 4641 25881 4675
rect 25881 4641 25915 4675
rect 25915 4641 25924 4675
rect 25872 4632 25924 4641
rect 26424 4675 26476 4684
rect 26424 4641 26433 4675
rect 26433 4641 26467 4675
rect 26467 4641 26476 4675
rect 26424 4632 26476 4641
rect 30748 4675 30800 4684
rect 30748 4641 30757 4675
rect 30757 4641 30791 4675
rect 30791 4641 30800 4675
rect 30748 4632 30800 4641
rect 36084 4675 36136 4684
rect 36084 4641 36093 4675
rect 36093 4641 36127 4675
rect 36127 4641 36136 4675
rect 36084 4632 36136 4641
rect 21456 4564 21508 4616
rect 22560 4564 22612 4616
rect 24124 4564 24176 4616
rect 28540 4607 28592 4616
rect 28540 4573 28549 4607
rect 28549 4573 28583 4607
rect 28583 4573 28592 4607
rect 28540 4564 28592 4573
rect 29000 4607 29052 4616
rect 29000 4573 29009 4607
rect 29009 4573 29043 4607
rect 29043 4573 29052 4607
rect 29000 4564 29052 4573
rect 34520 4564 34572 4616
rect 36728 4607 36780 4616
rect 36728 4573 36737 4607
rect 36737 4573 36771 4607
rect 36771 4573 36780 4607
rect 36728 4564 36780 4573
rect 34152 4496 34204 4548
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 24124 4088 24176 4140
rect 27436 4224 27488 4276
rect 25504 4088 25556 4140
rect 26148 4088 26200 4140
rect 28540 4088 28592 4140
rect 31300 4131 31352 4140
rect 31300 4097 31309 4131
rect 31309 4097 31343 4131
rect 31343 4097 31352 4131
rect 31300 4088 31352 4097
rect 34520 4131 34572 4140
rect 34520 4097 34529 4131
rect 34529 4097 34563 4131
rect 34563 4097 34572 4131
rect 34520 4088 34572 4097
rect 25872 4020 25924 4072
rect 26608 4063 26660 4072
rect 23664 3952 23716 4004
rect 26608 4029 26617 4063
rect 26617 4029 26651 4063
rect 26651 4029 26660 4063
rect 26608 4020 26660 4029
rect 29736 4063 29788 4072
rect 28908 3952 28960 4004
rect 19984 3884 20036 3936
rect 20628 3884 20680 3936
rect 22008 3884 22060 3936
rect 24492 3884 24544 3936
rect 24676 3927 24728 3936
rect 24676 3893 24685 3927
rect 24685 3893 24719 3927
rect 24719 3893 24728 3927
rect 24676 3884 24728 3893
rect 25412 3927 25464 3936
rect 25412 3893 25421 3927
rect 25421 3893 25455 3927
rect 25455 3893 25464 3927
rect 25412 3884 25464 3893
rect 26056 3927 26108 3936
rect 26056 3893 26065 3927
rect 26065 3893 26099 3927
rect 26099 3893 26108 3927
rect 26056 3884 26108 3893
rect 26148 3884 26200 3936
rect 26332 3884 26384 3936
rect 26516 3884 26568 3936
rect 29736 4029 29745 4063
rect 29745 4029 29779 4063
rect 29779 4029 29788 4063
rect 29736 4020 29788 4029
rect 33048 4063 33100 4072
rect 33048 4029 33057 4063
rect 33057 4029 33091 4063
rect 33091 4029 33100 4063
rect 33048 4020 33100 4029
rect 36728 4088 36780 4140
rect 30472 3952 30524 4004
rect 37188 3952 37240 4004
rect 31484 3884 31536 3936
rect 33416 3884 33468 3936
rect 35716 3884 35768 3936
rect 37280 3927 37332 3936
rect 37280 3893 37289 3927
rect 37289 3893 37323 3927
rect 37323 3893 37332 3927
rect 37280 3884 37332 3893
rect 38568 3884 38620 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 22836 3680 22888 3732
rect 26608 3680 26660 3732
rect 30840 3723 30892 3732
rect 30840 3689 30849 3723
rect 30849 3689 30883 3723
rect 30883 3689 30892 3723
rect 30840 3680 30892 3689
rect 36084 3680 36136 3732
rect 22284 3612 22336 3664
rect 9312 3476 9364 3528
rect 10784 3476 10836 3528
rect 12440 3476 12492 3528
rect 13544 3476 13596 3528
rect 14648 3476 14700 3528
rect 15476 3476 15528 3528
rect 16580 3476 16632 3528
rect 17316 3476 17368 3528
rect 18144 3476 18196 3528
rect 18972 3519 19024 3528
rect 18972 3485 18981 3519
rect 18981 3485 19015 3519
rect 19015 3485 19024 3519
rect 18972 3476 19024 3485
rect 20352 3476 20404 3528
rect 20904 3476 20956 3528
rect 22192 3476 22244 3528
rect 24124 3612 24176 3664
rect 24492 3612 24544 3664
rect 25320 3612 25372 3664
rect 25412 3612 25464 3664
rect 28356 3612 28408 3664
rect 36544 3612 36596 3664
rect 39948 3612 40000 3664
rect 29000 3544 29052 3596
rect 31484 3587 31536 3596
rect 23572 3519 23624 3528
rect 23572 3485 23581 3519
rect 23581 3485 23615 3519
rect 23615 3485 23624 3519
rect 23572 3476 23624 3485
rect 25872 3519 25924 3528
rect 25872 3485 25881 3519
rect 25881 3485 25915 3519
rect 25915 3485 25924 3519
rect 25872 3476 25924 3485
rect 27252 3476 27304 3528
rect 31484 3553 31493 3587
rect 31493 3553 31527 3587
rect 31527 3553 31536 3587
rect 31484 3544 31536 3553
rect 31944 3587 31996 3596
rect 31944 3553 31953 3587
rect 31953 3553 31987 3587
rect 31987 3553 31996 3587
rect 31944 3544 31996 3553
rect 34428 3587 34480 3596
rect 34428 3553 34437 3587
rect 34437 3553 34471 3587
rect 34471 3553 34480 3587
rect 34428 3544 34480 3553
rect 37280 3544 37332 3596
rect 37556 3544 37608 3596
rect 40776 3544 40828 3596
rect 36728 3519 36780 3528
rect 36728 3485 36737 3519
rect 36737 3485 36771 3519
rect 36771 3485 36780 3519
rect 36728 3476 36780 3485
rect 36820 3476 36872 3528
rect 39396 3476 39448 3528
rect 41328 3476 41380 3528
rect 42432 3476 42484 3528
rect 43260 3476 43312 3528
rect 44088 3476 44140 3528
rect 46020 3476 46072 3528
rect 46572 3476 46624 3528
rect 48228 3476 48280 3528
rect 49332 3476 49384 3528
rect 50160 3476 50212 3528
rect 52092 3476 52144 3528
rect 24308 3340 24360 3392
rect 26056 3340 26108 3392
rect 26516 3340 26568 3392
rect 26700 3408 26752 3460
rect 27804 3408 27856 3460
rect 29184 3408 29236 3460
rect 30656 3408 30708 3460
rect 37464 3408 37516 3460
rect 26976 3340 27028 3392
rect 33232 3340 33284 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 24676 3136 24728 3188
rect 30656 3179 30708 3188
rect 30656 3145 30665 3179
rect 30665 3145 30699 3179
rect 30699 3145 30708 3179
rect 30656 3136 30708 3145
rect 33232 3111 33284 3120
rect 33232 3077 33241 3111
rect 33241 3077 33275 3111
rect 33275 3077 33284 3111
rect 33232 3068 33284 3077
rect 16856 2932 16908 2984
rect 21180 2932 21232 2984
rect 22192 3043 22244 3052
rect 22192 3009 22201 3043
rect 22201 3009 22235 3043
rect 22235 3009 22244 3043
rect 22836 3043 22888 3052
rect 22192 3000 22244 3009
rect 22836 3009 22845 3043
rect 22845 3009 22879 3043
rect 22879 3009 22888 3043
rect 22836 3000 22888 3009
rect 24216 3000 24268 3052
rect 25504 3000 25556 3052
rect 23388 2932 23440 2984
rect 24676 2975 24728 2984
rect 24676 2941 24685 2975
rect 24685 2941 24719 2975
rect 24719 2941 24728 2975
rect 24676 2932 24728 2941
rect 25596 2975 25648 2984
rect 25596 2941 25605 2975
rect 25605 2941 25639 2975
rect 25639 2941 25648 2975
rect 25596 2932 25648 2941
rect 21732 2864 21784 2916
rect 24032 2864 24084 2916
rect 27620 3000 27672 3052
rect 27896 3043 27948 3052
rect 27896 3009 27905 3043
rect 27905 3009 27939 3043
rect 27939 3009 27948 3043
rect 27896 3000 27948 3009
rect 30472 3000 30524 3052
rect 31392 3000 31444 3052
rect 31760 3000 31812 3052
rect 33416 3043 33468 3052
rect 33416 3009 33425 3043
rect 33425 3009 33459 3043
rect 33459 3009 33468 3043
rect 33416 3000 33468 3009
rect 35716 3043 35768 3052
rect 35716 3009 35725 3043
rect 35725 3009 35759 3043
rect 35759 3009 35768 3043
rect 35716 3000 35768 3009
rect 36728 3000 36780 3052
rect 38016 3000 38068 3052
rect 40224 3000 40276 3052
rect 28632 2975 28684 2984
rect 7656 2796 7708 2848
rect 8576 2796 8628 2848
rect 9956 2796 10008 2848
rect 10508 2796 10560 2848
rect 11060 2796 11112 2848
rect 11612 2796 11664 2848
rect 12164 2839 12216 2848
rect 12164 2805 12173 2839
rect 12173 2805 12207 2839
rect 12207 2805 12216 2839
rect 12164 2796 12216 2805
rect 12992 2796 13044 2848
rect 13820 2796 13872 2848
rect 14372 2796 14424 2848
rect 15200 2796 15252 2848
rect 16028 2796 16080 2848
rect 17132 2796 17184 2848
rect 17868 2796 17920 2848
rect 18696 2796 18748 2848
rect 19432 2796 19484 2848
rect 25504 2796 25556 2848
rect 28632 2941 28641 2975
rect 28641 2941 28675 2975
rect 28675 2941 28684 2975
rect 28632 2932 28684 2941
rect 32220 2975 32272 2984
rect 32220 2941 32229 2975
rect 32229 2941 32263 2975
rect 32263 2941 32272 2975
rect 32220 2932 32272 2941
rect 33324 2864 33376 2916
rect 35348 2932 35400 2984
rect 39672 2932 39724 2984
rect 45468 2932 45520 2984
rect 46848 2932 46900 2984
rect 35808 2864 35860 2916
rect 38844 2864 38896 2916
rect 41052 2864 41104 2916
rect 42984 2864 43036 2916
rect 44364 2864 44416 2916
rect 47676 2864 47728 2916
rect 49056 2864 49108 2916
rect 50988 2864 51040 2916
rect 52368 2864 52420 2916
rect 29184 2796 29236 2848
rect 30012 2796 30064 2848
rect 30380 2796 30432 2848
rect 32772 2796 32824 2848
rect 34060 2796 34112 2848
rect 36176 2839 36228 2848
rect 36176 2805 36185 2839
rect 36185 2805 36219 2839
rect 36219 2805 36228 2839
rect 36176 2796 36228 2805
rect 36912 2796 36964 2848
rect 41880 2796 41932 2848
rect 43536 2796 43588 2848
rect 44916 2796 44968 2848
rect 46296 2796 46348 2848
rect 48504 2796 48556 2848
rect 49608 2796 49660 2848
rect 50620 2796 50672 2848
rect 51540 2796 51592 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 23572 2592 23624 2644
rect 25596 2592 25648 2644
rect 37464 2635 37516 2644
rect 37464 2601 37473 2635
rect 37473 2601 37507 2635
rect 37507 2601 37516 2635
rect 37464 2592 37516 2601
rect 38660 2635 38712 2644
rect 38660 2601 38669 2635
rect 38669 2601 38703 2635
rect 38703 2601 38712 2635
rect 38660 2592 38712 2601
rect 47952 2592 48004 2644
rect 9680 2524 9732 2576
rect 11336 2524 11388 2576
rect 14924 2524 14976 2576
rect 18420 2524 18472 2576
rect 20076 2524 20128 2576
rect 25044 2524 25096 2576
rect 34980 2524 35032 2576
rect 38292 2524 38344 2576
rect 41604 2524 41656 2576
rect 45192 2524 45244 2576
rect 48780 2524 48832 2576
rect 50712 2524 50764 2576
rect 12716 2456 12768 2508
rect 17592 2456 17644 2508
rect 19248 2456 19300 2508
rect 22836 2456 22888 2508
rect 27620 2456 27672 2508
rect 29460 2499 29512 2508
rect 29460 2465 29469 2499
rect 29469 2465 29503 2499
rect 29503 2465 29512 2499
rect 29460 2456 29512 2465
rect 31116 2499 31168 2508
rect 31116 2465 31125 2499
rect 31125 2465 31159 2499
rect 31159 2465 31168 2499
rect 31116 2456 31168 2465
rect 31760 2456 31812 2508
rect 36176 2456 36228 2508
rect 39120 2456 39172 2508
rect 8208 2388 8260 2440
rect 8944 2388 8996 2440
rect 10232 2388 10284 2440
rect 11888 2388 11940 2440
rect 13268 2388 13320 2440
rect 14096 2388 14148 2440
rect 16304 2388 16356 2440
rect 15752 2320 15804 2372
rect 24124 2388 24176 2440
rect 24216 2431 24268 2440
rect 24216 2397 24225 2431
rect 24225 2397 24259 2431
rect 24259 2397 24268 2431
rect 24216 2388 24268 2397
rect 36544 2388 36596 2440
rect 36728 2388 36780 2440
rect 42156 2456 42208 2508
rect 44640 2456 44692 2508
rect 47124 2456 47176 2508
rect 49884 2456 49936 2508
rect 51816 2456 51868 2508
rect 23756 2320 23808 2372
rect 24032 2320 24084 2372
rect 27252 2320 27304 2372
rect 33600 2320 33652 2372
rect 36360 2252 36412 2304
rect 37740 2320 37792 2372
rect 40500 2320 40552 2372
rect 42708 2388 42760 2440
rect 43812 2320 43864 2372
rect 45744 2388 45796 2440
rect 47400 2320 47452 2372
rect 51264 2320 51316 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 24124 2048 24176 2100
rect 25872 2048 25924 2100
rect 23756 1368 23808 1420
rect 24492 1368 24544 1420
<< metal2 >>
rect 3698 59200 3754 60000
rect 4158 59200 4214 60000
rect 4618 59200 4674 60000
rect 5078 59200 5134 60000
rect 5538 59200 5594 60000
rect 5998 59200 6054 60000
rect 6458 59200 6514 60000
rect 6918 59200 6974 60000
rect 7378 59200 7434 60000
rect 7838 59200 7894 60000
rect 8298 59200 8354 60000
rect 8758 59200 8814 60000
rect 9218 59200 9274 60000
rect 9678 59200 9734 60000
rect 10138 59200 10194 60000
rect 10598 59200 10654 60000
rect 11058 59200 11114 60000
rect 11518 59200 11574 60000
rect 11978 59200 12034 60000
rect 12438 59200 12494 60000
rect 12898 59200 12954 60000
rect 13358 59200 13414 60000
rect 13818 59200 13874 60000
rect 14278 59200 14334 60000
rect 14738 59200 14794 60000
rect 15198 59200 15254 60000
rect 15658 59200 15714 60000
rect 16118 59200 16174 60000
rect 16578 59200 16634 60000
rect 17038 59200 17094 60000
rect 17498 59200 17554 60000
rect 17958 59200 18014 60000
rect 18418 59200 18474 60000
rect 18878 59200 18934 60000
rect 19338 59200 19394 60000
rect 19798 59200 19854 60000
rect 20258 59200 20314 60000
rect 20718 59200 20774 60000
rect 21178 59200 21234 60000
rect 21638 59200 21694 60000
rect 21744 59214 22048 59242
rect 3712 57594 3740 59200
rect 3700 57588 3752 57594
rect 3700 57530 3752 57536
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4632 57050 4660 59200
rect 5092 57594 5120 59200
rect 5080 57588 5132 57594
rect 5080 57530 5132 57536
rect 6012 57458 6040 59200
rect 6472 57458 6500 59200
rect 7392 57458 7420 59200
rect 7852 57458 7880 59200
rect 8772 57458 8800 59200
rect 9232 57458 9260 59200
rect 5448 57452 5500 57458
rect 5448 57394 5500 57400
rect 6000 57452 6052 57458
rect 6000 57394 6052 57400
rect 6460 57452 6512 57458
rect 6460 57394 6512 57400
rect 7380 57452 7432 57458
rect 7380 57394 7432 57400
rect 7840 57452 7892 57458
rect 7840 57394 7892 57400
rect 8760 57452 8812 57458
rect 8760 57394 8812 57400
rect 9220 57452 9272 57458
rect 9220 57394 9272 57400
rect 5356 57316 5408 57322
rect 5356 57258 5408 57264
rect 4620 57044 4672 57050
rect 4620 56986 4672 56992
rect 5368 56166 5396 57258
rect 5460 56710 5488 57394
rect 10152 57050 10180 59200
rect 10612 57594 10640 59200
rect 10600 57588 10652 57594
rect 10600 57530 10652 57536
rect 11532 57458 11560 59200
rect 11992 57594 12020 59200
rect 12348 57860 12400 57866
rect 12348 57802 12400 57808
rect 11980 57588 12032 57594
rect 11980 57530 12032 57536
rect 12360 57458 12388 57802
rect 10968 57452 11020 57458
rect 10968 57394 11020 57400
rect 11520 57452 11572 57458
rect 11520 57394 11572 57400
rect 12348 57452 12400 57458
rect 12348 57394 12400 57400
rect 10140 57044 10192 57050
rect 10140 56986 10192 56992
rect 10980 56982 11008 57394
rect 12912 57050 12940 59200
rect 13372 57594 13400 59200
rect 13360 57588 13412 57594
rect 13360 57530 13412 57536
rect 14292 57458 14320 59200
rect 14752 57594 14780 59200
rect 15108 57928 15160 57934
rect 15108 57870 15160 57876
rect 14740 57588 14792 57594
rect 14740 57530 14792 57536
rect 15120 57458 15148 57870
rect 14280 57452 14332 57458
rect 14280 57394 14332 57400
rect 15108 57452 15160 57458
rect 15108 57394 15160 57400
rect 15672 57050 15700 59200
rect 16132 57594 16160 59200
rect 16120 57588 16172 57594
rect 16120 57530 16172 57536
rect 17052 57458 17080 59200
rect 17512 57594 17540 59200
rect 17500 57588 17552 57594
rect 17500 57530 17552 57536
rect 18432 57458 18460 59200
rect 18892 57594 18920 59200
rect 19812 58018 19840 59200
rect 19812 57990 20024 58018
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 18880 57588 18932 57594
rect 18880 57530 18932 57536
rect 16488 57452 16540 57458
rect 16488 57394 16540 57400
rect 17040 57452 17092 57458
rect 17040 57394 17092 57400
rect 17868 57452 17920 57458
rect 17868 57394 17920 57400
rect 18420 57452 18472 57458
rect 18420 57394 18472 57400
rect 12900 57044 12952 57050
rect 12900 56986 12952 56992
rect 15660 57044 15712 57050
rect 15660 56986 15712 56992
rect 10968 56976 11020 56982
rect 10968 56918 11020 56924
rect 16500 56914 16528 57394
rect 16488 56908 16540 56914
rect 16488 56850 16540 56856
rect 5448 56704 5500 56710
rect 5448 56646 5500 56652
rect 17880 56438 17908 57394
rect 19996 57050 20024 57990
rect 20272 57594 20300 59200
rect 20260 57588 20312 57594
rect 20260 57530 20312 57536
rect 20628 57452 20680 57458
rect 20628 57394 20680 57400
rect 20640 57254 20668 57394
rect 20628 57248 20680 57254
rect 20628 57190 20680 57196
rect 21192 57050 21220 59200
rect 21652 59106 21680 59200
rect 21744 59106 21772 59214
rect 21652 59078 21772 59106
rect 22020 57576 22048 59214
rect 22098 59200 22154 60000
rect 22558 59200 22614 60000
rect 23018 59200 23074 60000
rect 23478 59200 23534 60000
rect 23938 59200 23994 60000
rect 24398 59200 24454 60000
rect 24504 59214 24808 59242
rect 22100 57588 22152 57594
rect 22020 57548 22100 57576
rect 22100 57530 22152 57536
rect 21454 57488 21510 57497
rect 21454 57423 21510 57432
rect 22284 57452 22336 57458
rect 21468 57322 21496 57423
rect 22284 57394 22336 57400
rect 21456 57316 21508 57322
rect 21456 57258 21508 57264
rect 19984 57044 20036 57050
rect 19984 56986 20036 56992
rect 21180 57044 21232 57050
rect 21180 56986 21232 56992
rect 22296 56681 22324 57394
rect 22282 56672 22338 56681
rect 19574 56604 19882 56613
rect 22282 56607 22338 56616
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 17868 56432 17920 56438
rect 17868 56374 17920 56380
rect 22572 56370 22600 59200
rect 23032 57594 23060 59200
rect 23204 57996 23256 58002
rect 23204 57938 23256 57944
rect 23020 57588 23072 57594
rect 23020 57530 23072 57536
rect 23216 57050 23244 57938
rect 23756 57792 23808 57798
rect 23756 57734 23808 57740
rect 23388 57452 23440 57458
rect 23308 57412 23388 57440
rect 23204 57044 23256 57050
rect 23204 56986 23256 56992
rect 23308 56545 23336 57412
rect 23388 57394 23440 57400
rect 23388 57316 23440 57322
rect 23388 57258 23440 57264
rect 23400 56846 23428 57258
rect 23480 57044 23532 57050
rect 23480 56986 23532 56992
rect 23388 56840 23440 56846
rect 23388 56782 23440 56788
rect 23294 56536 23350 56545
rect 23294 56471 23350 56480
rect 22560 56364 22612 56370
rect 22560 56306 22612 56312
rect 5356 56160 5408 56166
rect 5356 56102 5408 56108
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 23400 55418 23428 56782
rect 23492 56506 23520 56986
rect 23768 56710 23796 57734
rect 23952 57497 23980 59200
rect 24412 59106 24440 59200
rect 24504 59106 24532 59214
rect 24412 59078 24532 59106
rect 24780 57576 24808 59214
rect 24858 59200 24914 60000
rect 25318 59200 25374 60000
rect 25778 59200 25834 60000
rect 26238 59200 26294 60000
rect 26698 59200 26754 60000
rect 27158 59200 27214 60000
rect 27618 59200 27674 60000
rect 28078 59200 28134 60000
rect 28538 59200 28594 60000
rect 28998 59200 29054 60000
rect 29458 59200 29514 60000
rect 29918 59200 29974 60000
rect 30378 59200 30434 60000
rect 30838 59200 30894 60000
rect 31298 59200 31354 60000
rect 31758 59200 31814 60000
rect 32218 59200 32274 60000
rect 32678 59200 32734 60000
rect 33138 59200 33194 60000
rect 33598 59200 33654 60000
rect 34058 59200 34114 60000
rect 34518 59200 34574 60000
rect 34978 59200 35034 60000
rect 35084 59214 35388 59242
rect 25044 57928 25096 57934
rect 25044 57870 25096 57876
rect 24860 57588 24912 57594
rect 24780 57548 24860 57576
rect 24860 57530 24912 57536
rect 23938 57488 23994 57497
rect 23938 57423 23994 57432
rect 24032 57452 24084 57458
rect 24032 57394 24084 57400
rect 24124 57452 24176 57458
rect 24124 57394 24176 57400
rect 23940 57384 23992 57390
rect 23940 57326 23992 57332
rect 23848 57248 23900 57254
rect 23848 57190 23900 57196
rect 23756 56704 23808 56710
rect 23756 56646 23808 56652
rect 23480 56500 23532 56506
rect 23480 56442 23532 56448
rect 23768 55758 23796 56646
rect 23860 56370 23888 57190
rect 23952 56710 23980 57326
rect 24044 56846 24072 57394
rect 24136 57050 24164 57394
rect 24308 57384 24360 57390
rect 24308 57326 24360 57332
rect 24584 57384 24636 57390
rect 24584 57326 24636 57332
rect 24124 57044 24176 57050
rect 24124 56986 24176 56992
rect 24032 56840 24084 56846
rect 24032 56782 24084 56788
rect 23940 56704 23992 56710
rect 23940 56646 23992 56652
rect 23848 56364 23900 56370
rect 23848 56306 23900 56312
rect 24320 56302 24348 57326
rect 24596 57050 24624 57326
rect 25056 57050 25084 57870
rect 24584 57044 24636 57050
rect 24584 56986 24636 56992
rect 25044 57044 25096 57050
rect 25044 56986 25096 56992
rect 25332 56982 25360 59200
rect 25792 57594 25820 59200
rect 25780 57588 25832 57594
rect 25780 57530 25832 57536
rect 25596 57452 25648 57458
rect 25596 57394 25648 57400
rect 25320 56976 25372 56982
rect 25320 56918 25372 56924
rect 25608 56846 25636 57394
rect 26332 57384 26384 57390
rect 26332 57326 26384 57332
rect 25688 57248 25740 57254
rect 25688 57190 25740 57196
rect 25700 56846 25728 57190
rect 25412 56840 25464 56846
rect 25412 56782 25464 56788
rect 25596 56840 25648 56846
rect 25596 56782 25648 56788
rect 25688 56840 25740 56846
rect 25688 56782 25740 56788
rect 24308 56296 24360 56302
rect 24308 56238 24360 56244
rect 24768 56296 24820 56302
rect 24768 56238 24820 56244
rect 24780 55826 24808 56238
rect 24768 55820 24820 55826
rect 24768 55762 24820 55768
rect 23756 55752 23808 55758
rect 23756 55694 23808 55700
rect 24032 55616 24084 55622
rect 24032 55558 24084 55564
rect 23388 55412 23440 55418
rect 23388 55354 23440 55360
rect 24044 55282 24072 55558
rect 24032 55276 24084 55282
rect 24032 55218 24084 55224
rect 24780 55078 24808 55762
rect 25424 55758 25452 56782
rect 25504 56704 25556 56710
rect 25504 56646 25556 56652
rect 25516 56409 25544 56646
rect 25502 56400 25558 56409
rect 25502 56335 25504 56344
rect 25556 56335 25558 56344
rect 25504 56306 25556 56312
rect 25608 55962 25636 56782
rect 25700 56250 25728 56782
rect 26238 56672 26294 56681
rect 26238 56607 26294 56616
rect 26252 56370 26280 56607
rect 26240 56364 26292 56370
rect 26240 56306 26292 56312
rect 25700 56222 25820 56250
rect 25688 56160 25740 56166
rect 25688 56102 25740 56108
rect 25596 55956 25648 55962
rect 25596 55898 25648 55904
rect 25412 55752 25464 55758
rect 25412 55694 25464 55700
rect 25700 55282 25728 56102
rect 25792 55418 25820 56222
rect 26252 55418 26280 56306
rect 26344 56234 26372 57326
rect 26516 56840 26568 56846
rect 26516 56782 26568 56788
rect 26608 56840 26660 56846
rect 26608 56782 26660 56788
rect 26424 56704 26476 56710
rect 26424 56646 26476 56652
rect 26332 56228 26384 56234
rect 26332 56170 26384 56176
rect 26344 55962 26372 56170
rect 26332 55956 26384 55962
rect 26332 55898 26384 55904
rect 25780 55412 25832 55418
rect 25780 55354 25832 55360
rect 26240 55412 26292 55418
rect 26240 55354 26292 55360
rect 26436 55282 26464 56646
rect 26528 56506 26556 56782
rect 26516 56500 26568 56506
rect 26516 56442 26568 56448
rect 26620 56166 26648 56782
rect 26608 56160 26660 56166
rect 26608 56102 26660 56108
rect 26620 55282 26648 56102
rect 25688 55276 25740 55282
rect 25688 55218 25740 55224
rect 26424 55276 26476 55282
rect 26424 55218 26476 55224
rect 26608 55276 26660 55282
rect 26608 55218 26660 55224
rect 24768 55072 24820 55078
rect 24768 55014 24820 55020
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 24780 54806 24808 55014
rect 26620 54874 26648 55218
rect 26712 54874 26740 59200
rect 26976 57860 27028 57866
rect 26976 57802 27028 57808
rect 27068 57860 27120 57866
rect 27068 57802 27120 57808
rect 26988 56914 27016 57802
rect 26884 56908 26936 56914
rect 26884 56850 26936 56856
rect 26976 56908 27028 56914
rect 26976 56850 27028 56856
rect 26896 56506 26924 56850
rect 27080 56846 27108 57802
rect 27172 57594 27200 59200
rect 27160 57588 27212 57594
rect 27160 57530 27212 57536
rect 27160 57452 27212 57458
rect 27160 57394 27212 57400
rect 27804 57452 27856 57458
rect 27804 57394 27856 57400
rect 27172 57338 27200 57394
rect 27172 57310 27568 57338
rect 27172 57254 27200 57310
rect 27540 57254 27568 57310
rect 27160 57248 27212 57254
rect 27160 57190 27212 57196
rect 27436 57248 27488 57254
rect 27436 57190 27488 57196
rect 27528 57248 27580 57254
rect 27528 57190 27580 57196
rect 27068 56840 27120 56846
rect 27068 56782 27120 56788
rect 26884 56500 26936 56506
rect 26884 56442 26936 56448
rect 26976 56432 27028 56438
rect 26976 56374 27028 56380
rect 26884 56364 26936 56370
rect 26884 56306 26936 56312
rect 26896 55894 26924 56306
rect 26884 55888 26936 55894
rect 26988 55865 27016 56374
rect 26884 55830 26936 55836
rect 26974 55856 27030 55865
rect 26974 55791 27030 55800
rect 26976 55752 27028 55758
rect 26976 55694 27028 55700
rect 26608 54868 26660 54874
rect 26608 54810 26660 54816
rect 26700 54868 26752 54874
rect 26700 54810 26752 54816
rect 26988 54806 27016 55694
rect 24768 54800 24820 54806
rect 24768 54742 24820 54748
rect 26976 54800 27028 54806
rect 26976 54742 27028 54748
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 26988 54058 27016 54742
rect 27080 54330 27108 56782
rect 27344 56704 27396 56710
rect 27344 56646 27396 56652
rect 27356 56370 27384 56646
rect 27448 56438 27476 57190
rect 27816 57050 27844 57394
rect 27804 57044 27856 57050
rect 27804 56986 27856 56992
rect 27528 56840 27580 56846
rect 27528 56782 27580 56788
rect 27712 56840 27764 56846
rect 27712 56782 27764 56788
rect 27436 56432 27488 56438
rect 27436 56374 27488 56380
rect 27344 56364 27396 56370
rect 27344 56306 27396 56312
rect 27540 55706 27568 56782
rect 27724 56506 27752 56782
rect 27712 56500 27764 56506
rect 27712 56442 27764 56448
rect 27620 56364 27672 56370
rect 27620 56306 27672 56312
rect 27712 56364 27764 56370
rect 27712 56306 27764 56312
rect 27632 56166 27660 56306
rect 27620 56160 27672 56166
rect 27620 56102 27672 56108
rect 27540 55678 27660 55706
rect 27528 55276 27580 55282
rect 27528 55218 27580 55224
rect 27068 54324 27120 54330
rect 27068 54266 27120 54272
rect 26976 54052 27028 54058
rect 26976 53994 27028 54000
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 27540 52426 27568 55218
rect 27632 55078 27660 55678
rect 27724 55282 27752 56306
rect 27896 55684 27948 55690
rect 27896 55626 27948 55632
rect 27712 55276 27764 55282
rect 27712 55218 27764 55224
rect 27620 55072 27672 55078
rect 27620 55014 27672 55020
rect 27908 54330 27936 55626
rect 28092 54874 28120 59200
rect 28552 57594 28580 59200
rect 28540 57588 28592 57594
rect 28540 57530 28592 57536
rect 28816 57248 28868 57254
rect 28816 57190 28868 57196
rect 28172 56976 28224 56982
rect 28172 56918 28224 56924
rect 28184 56370 28212 56918
rect 28828 56846 28856 57190
rect 28908 56976 28960 56982
rect 28908 56918 28960 56924
rect 28724 56840 28776 56846
rect 28724 56782 28776 56788
rect 28816 56840 28868 56846
rect 28816 56782 28868 56788
rect 28356 56772 28408 56778
rect 28356 56714 28408 56720
rect 28264 56500 28316 56506
rect 28264 56442 28316 56448
rect 28172 56364 28224 56370
rect 28172 56306 28224 56312
rect 28276 55826 28304 56442
rect 28264 55820 28316 55826
rect 28264 55762 28316 55768
rect 28368 55418 28396 56714
rect 28540 56704 28592 56710
rect 28540 56646 28592 56652
rect 28448 56364 28500 56370
rect 28448 56306 28500 56312
rect 28460 55826 28488 56306
rect 28552 55826 28580 56646
rect 28448 55820 28500 55826
rect 28448 55762 28500 55768
rect 28540 55820 28592 55826
rect 28540 55762 28592 55768
rect 28356 55412 28408 55418
rect 28356 55354 28408 55360
rect 28460 55282 28488 55762
rect 28448 55276 28500 55282
rect 28448 55218 28500 55224
rect 28552 55214 28580 55762
rect 28632 55752 28684 55758
rect 28736 55706 28764 56782
rect 28684 55700 28764 55706
rect 28632 55694 28764 55700
rect 28816 55752 28868 55758
rect 28816 55694 28868 55700
rect 28644 55678 28764 55694
rect 28540 55208 28592 55214
rect 28540 55150 28592 55156
rect 28448 55072 28500 55078
rect 28448 55014 28500 55020
rect 28080 54868 28132 54874
rect 28080 54810 28132 54816
rect 27896 54324 27948 54330
rect 27896 54266 27948 54272
rect 28460 54126 28488 55014
rect 28736 54874 28764 55678
rect 28828 55418 28856 55694
rect 28816 55412 28868 55418
rect 28816 55354 28868 55360
rect 28724 54868 28776 54874
rect 28724 54810 28776 54816
rect 28540 54800 28592 54806
rect 28540 54742 28592 54748
rect 28552 54194 28580 54742
rect 28920 54330 28948 56918
rect 29012 55690 29040 59200
rect 29092 57452 29144 57458
rect 29092 57394 29144 57400
rect 29104 57050 29132 57394
rect 29184 57316 29236 57322
rect 29184 57258 29236 57264
rect 29196 57050 29224 57258
rect 29092 57044 29144 57050
rect 29092 56986 29144 56992
rect 29184 57044 29236 57050
rect 29184 56986 29236 56992
rect 29104 56352 29132 56986
rect 29184 56908 29236 56914
rect 29184 56850 29236 56856
rect 29196 56710 29224 56850
rect 29276 56840 29328 56846
rect 29274 56808 29276 56817
rect 29328 56808 29330 56817
rect 29330 56766 29408 56794
rect 29274 56743 29330 56752
rect 29184 56704 29236 56710
rect 29184 56646 29236 56652
rect 29274 56536 29330 56545
rect 29274 56471 29330 56480
rect 29288 56438 29316 56471
rect 29276 56432 29328 56438
rect 29276 56374 29328 56380
rect 29184 56364 29236 56370
rect 29104 56324 29184 56352
rect 29184 56306 29236 56312
rect 29380 55826 29408 56766
rect 29368 55820 29420 55826
rect 29368 55762 29420 55768
rect 29472 55706 29500 59200
rect 29552 57520 29604 57526
rect 29552 57462 29604 57468
rect 29564 56914 29592 57462
rect 29552 56908 29604 56914
rect 29552 56850 29604 56856
rect 29564 56166 29592 56850
rect 29828 56840 29880 56846
rect 29828 56782 29880 56788
rect 29840 56506 29868 56782
rect 29828 56500 29880 56506
rect 29828 56442 29880 56448
rect 29932 56370 29960 59200
rect 30392 57458 30420 59200
rect 30852 57458 30880 59200
rect 30380 57452 30432 57458
rect 30380 57394 30432 57400
rect 30840 57452 30892 57458
rect 30840 57394 30892 57400
rect 31312 57390 31340 59200
rect 31772 57458 31800 59200
rect 31760 57452 31812 57458
rect 31760 57394 31812 57400
rect 31300 57384 31352 57390
rect 31300 57326 31352 57332
rect 30656 56908 30708 56914
rect 30656 56850 30708 56856
rect 31116 56908 31168 56914
rect 31116 56850 31168 56856
rect 30668 56817 30696 56850
rect 30932 56840 30984 56846
rect 30654 56808 30710 56817
rect 30932 56782 30984 56788
rect 30654 56743 30710 56752
rect 30104 56432 30156 56438
rect 30104 56374 30156 56380
rect 29920 56364 29972 56370
rect 29920 56306 29972 56312
rect 29552 56160 29604 56166
rect 29552 56102 29604 56108
rect 29920 55820 29972 55826
rect 29920 55762 29972 55768
rect 29736 55752 29788 55758
rect 29000 55684 29052 55690
rect 29472 55678 29592 55706
rect 29736 55694 29788 55700
rect 29000 55626 29052 55632
rect 29276 55616 29328 55622
rect 29274 55584 29276 55593
rect 29460 55616 29512 55622
rect 29328 55584 29330 55593
rect 29460 55558 29512 55564
rect 29274 55519 29330 55528
rect 29472 55350 29500 55558
rect 29460 55344 29512 55350
rect 29460 55286 29512 55292
rect 29184 54596 29236 54602
rect 29184 54538 29236 54544
rect 29000 54528 29052 54534
rect 29000 54470 29052 54476
rect 28908 54324 28960 54330
rect 28908 54266 28960 54272
rect 28540 54188 28592 54194
rect 28540 54130 28592 54136
rect 28448 54120 28500 54126
rect 28448 54062 28500 54068
rect 28632 54052 28684 54058
rect 28632 53994 28684 54000
rect 28644 53446 28672 53994
rect 29012 53786 29040 54470
rect 29196 54330 29224 54538
rect 29472 54534 29500 55286
rect 29564 54874 29592 55678
rect 29748 55350 29776 55694
rect 29932 55350 29960 55762
rect 30116 55758 30144 56374
rect 30668 56166 30696 56743
rect 30944 56166 30972 56782
rect 31128 56302 31156 56850
rect 31208 56840 31260 56846
rect 31208 56782 31260 56788
rect 31220 56506 31248 56782
rect 31760 56704 31812 56710
rect 31760 56646 31812 56652
rect 31944 56704 31996 56710
rect 31944 56646 31996 56652
rect 31208 56500 31260 56506
rect 31208 56442 31260 56448
rect 31772 56370 31800 56646
rect 31760 56364 31812 56370
rect 31760 56306 31812 56312
rect 31116 56296 31168 56302
rect 31116 56238 31168 56244
rect 31576 56296 31628 56302
rect 31576 56238 31628 56244
rect 30656 56160 30708 56166
rect 30656 56102 30708 56108
rect 30932 56160 30984 56166
rect 30932 56102 30984 56108
rect 30104 55752 30156 55758
rect 30104 55694 30156 55700
rect 30668 55622 30696 56102
rect 30944 55962 30972 56102
rect 30932 55956 30984 55962
rect 30932 55898 30984 55904
rect 30840 55752 30892 55758
rect 30840 55694 30892 55700
rect 31300 55752 31352 55758
rect 31300 55694 31352 55700
rect 30748 55684 30800 55690
rect 30748 55626 30800 55632
rect 30656 55616 30708 55622
rect 30656 55558 30708 55564
rect 30760 55418 30788 55626
rect 30748 55412 30800 55418
rect 30748 55354 30800 55360
rect 29736 55344 29788 55350
rect 29736 55286 29788 55292
rect 29920 55344 29972 55350
rect 29920 55286 29972 55292
rect 30380 55276 30432 55282
rect 30380 55218 30432 55224
rect 30564 55276 30616 55282
rect 30564 55218 30616 55224
rect 29552 54868 29604 54874
rect 29552 54810 29604 54816
rect 30392 54806 30420 55218
rect 30380 54800 30432 54806
rect 30380 54742 30432 54748
rect 30392 54670 30420 54742
rect 29644 54664 29696 54670
rect 29644 54606 29696 54612
rect 30380 54664 30432 54670
rect 30380 54606 30432 54612
rect 29460 54528 29512 54534
rect 29460 54470 29512 54476
rect 29656 54330 29684 54606
rect 30576 54602 30604 55218
rect 30852 54874 30880 55694
rect 31116 55684 31168 55690
rect 31116 55626 31168 55632
rect 30840 54868 30892 54874
rect 30840 54810 30892 54816
rect 31128 54602 31156 55626
rect 31312 55418 31340 55694
rect 31300 55412 31352 55418
rect 31300 55354 31352 55360
rect 31588 55282 31616 56238
rect 31852 56160 31904 56166
rect 31956 56148 31984 56646
rect 32232 56370 32260 59200
rect 32404 57384 32456 57390
rect 32404 57326 32456 57332
rect 32312 56840 32364 56846
rect 32312 56782 32364 56788
rect 32220 56364 32272 56370
rect 32220 56306 32272 56312
rect 31904 56120 31984 56148
rect 31852 56102 31904 56108
rect 31576 55276 31628 55282
rect 31576 55218 31628 55224
rect 31864 55078 31892 56102
rect 32324 55622 32352 56782
rect 32416 55758 32444 57326
rect 32692 57050 32720 59200
rect 33152 57594 33180 59200
rect 33612 58018 33640 59200
rect 33612 57990 33824 58018
rect 33692 57860 33744 57866
rect 33692 57802 33744 57808
rect 33140 57588 33192 57594
rect 33140 57530 33192 57536
rect 32772 57452 32824 57458
rect 32772 57394 32824 57400
rect 33600 57452 33652 57458
rect 33600 57394 33652 57400
rect 32680 57044 32732 57050
rect 32680 56986 32732 56992
rect 32784 56846 32812 57394
rect 32956 57384 33008 57390
rect 32956 57326 33008 57332
rect 32772 56840 32824 56846
rect 32772 56782 32824 56788
rect 32968 56828 32996 57326
rect 33048 57248 33100 57254
rect 33324 57248 33376 57254
rect 33100 57208 33180 57236
rect 33048 57190 33100 57196
rect 33048 56840 33100 56846
rect 32968 56800 33048 56828
rect 32968 56438 32996 56800
rect 33048 56782 33100 56788
rect 32956 56432 33008 56438
rect 32956 56374 33008 56380
rect 33152 56302 33180 57208
rect 33324 57190 33376 57196
rect 33336 56982 33364 57190
rect 33324 56976 33376 56982
rect 33324 56918 33376 56924
rect 33336 56370 33364 56918
rect 33612 56370 33640 57394
rect 33704 56710 33732 57802
rect 33692 56704 33744 56710
rect 33692 56646 33744 56652
rect 33324 56364 33376 56370
rect 33324 56306 33376 56312
rect 33600 56364 33652 56370
rect 33600 56306 33652 56312
rect 33140 56296 33192 56302
rect 33140 56238 33192 56244
rect 33048 56160 33100 56166
rect 33048 56102 33100 56108
rect 33060 55758 33088 56102
rect 32404 55752 32456 55758
rect 32404 55694 32456 55700
rect 32680 55752 32732 55758
rect 32680 55694 32732 55700
rect 33048 55752 33100 55758
rect 33048 55694 33100 55700
rect 32312 55616 32364 55622
rect 32312 55558 32364 55564
rect 32324 55214 32352 55558
rect 32692 55282 32720 55694
rect 32864 55684 32916 55690
rect 32864 55626 32916 55632
rect 32876 55593 32904 55626
rect 32862 55584 32918 55593
rect 32862 55519 32918 55528
rect 32680 55276 32732 55282
rect 32680 55218 32732 55224
rect 32312 55208 32364 55214
rect 32312 55150 32364 55156
rect 31852 55072 31904 55078
rect 31852 55014 31904 55020
rect 32404 55072 32456 55078
rect 32404 55014 32456 55020
rect 32416 54670 32444 55014
rect 32404 54664 32456 54670
rect 32324 54612 32404 54618
rect 32324 54606 32456 54612
rect 30564 54596 30616 54602
rect 30564 54538 30616 54544
rect 31116 54596 31168 54602
rect 31116 54538 31168 54544
rect 32324 54590 32444 54606
rect 32588 54596 32640 54602
rect 29184 54324 29236 54330
rect 29184 54266 29236 54272
rect 29644 54324 29696 54330
rect 29644 54266 29696 54272
rect 29736 54256 29788 54262
rect 29736 54198 29788 54204
rect 29748 54126 29776 54198
rect 30576 54126 30604 54538
rect 29736 54120 29788 54126
rect 29736 54062 29788 54068
rect 30564 54120 30616 54126
rect 30564 54062 30616 54068
rect 29000 53780 29052 53786
rect 29000 53722 29052 53728
rect 29748 53582 29776 54062
rect 30196 54052 30248 54058
rect 30196 53994 30248 54000
rect 30208 53582 30236 53994
rect 31128 53990 31156 54538
rect 32324 54126 32352 54590
rect 32588 54538 32640 54544
rect 32404 54188 32456 54194
rect 32404 54130 32456 54136
rect 32312 54120 32364 54126
rect 32312 54062 32364 54068
rect 31116 53984 31168 53990
rect 31116 53926 31168 53932
rect 31128 53718 31156 53926
rect 32416 53786 32444 54130
rect 32600 53786 32628 54538
rect 32692 54262 32720 55218
rect 33152 54670 33180 56238
rect 33336 56166 33364 56306
rect 33324 56160 33376 56166
rect 33324 56102 33376 56108
rect 33232 55752 33284 55758
rect 33232 55694 33284 55700
rect 33140 54664 33192 54670
rect 33140 54606 33192 54612
rect 32864 54528 32916 54534
rect 32864 54470 32916 54476
rect 32680 54256 32732 54262
rect 32680 54198 32732 54204
rect 32404 53780 32456 53786
rect 32404 53722 32456 53728
rect 32588 53780 32640 53786
rect 32588 53722 32640 53728
rect 31116 53712 31168 53718
rect 31116 53654 31168 53660
rect 32876 53582 32904 54470
rect 33152 53650 33180 54606
rect 33244 54330 33272 55694
rect 33336 55282 33364 56102
rect 33612 55350 33640 56306
rect 33796 55962 33824 57990
rect 33784 55956 33836 55962
rect 33784 55898 33836 55904
rect 34072 55758 34100 59200
rect 34532 57458 34560 59200
rect 34992 59106 35020 59200
rect 35084 59106 35112 59214
rect 34992 59078 35112 59106
rect 34244 57452 34296 57458
rect 34244 57394 34296 57400
rect 34520 57452 34572 57458
rect 34520 57394 34572 57400
rect 34704 57452 34756 57458
rect 34704 57394 34756 57400
rect 34256 57254 34284 57394
rect 34336 57384 34388 57390
rect 34336 57326 34388 57332
rect 34612 57384 34664 57390
rect 34612 57326 34664 57332
rect 34244 57248 34296 57254
rect 34244 57190 34296 57196
rect 34348 56846 34376 57326
rect 34336 56840 34388 56846
rect 34336 56782 34388 56788
rect 34520 56840 34572 56846
rect 34520 56782 34572 56788
rect 33692 55752 33744 55758
rect 33692 55694 33744 55700
rect 34060 55752 34112 55758
rect 34060 55694 34112 55700
rect 33600 55344 33652 55350
rect 33600 55286 33652 55292
rect 33704 55282 33732 55694
rect 34348 55690 34376 56782
rect 34336 55684 34388 55690
rect 34336 55626 34388 55632
rect 34348 55350 34376 55626
rect 34336 55344 34388 55350
rect 34336 55286 34388 55292
rect 33324 55276 33376 55282
rect 33324 55218 33376 55224
rect 33692 55276 33744 55282
rect 33692 55218 33744 55224
rect 33324 54664 33376 54670
rect 33324 54606 33376 54612
rect 33336 54330 33364 54606
rect 33508 54528 33560 54534
rect 33508 54470 33560 54476
rect 33232 54324 33284 54330
rect 33232 54266 33284 54272
rect 33324 54324 33376 54330
rect 33324 54266 33376 54272
rect 33140 53644 33192 53650
rect 33140 53586 33192 53592
rect 33336 53582 33364 54266
rect 33520 53786 33548 54470
rect 33704 53990 33732 55218
rect 34428 55208 34480 55214
rect 34428 55150 34480 55156
rect 33876 54732 33928 54738
rect 33876 54674 33928 54680
rect 33888 54126 33916 54674
rect 34440 54670 34468 55150
rect 34428 54664 34480 54670
rect 34428 54606 34480 54612
rect 34440 54194 34468 54606
rect 34428 54188 34480 54194
rect 34428 54130 34480 54136
rect 33876 54120 33928 54126
rect 33876 54062 33928 54068
rect 33692 53984 33744 53990
rect 33692 53926 33744 53932
rect 33508 53780 33560 53786
rect 33508 53722 33560 53728
rect 33704 53718 33732 53926
rect 33692 53712 33744 53718
rect 33692 53654 33744 53660
rect 29736 53576 29788 53582
rect 29736 53518 29788 53524
rect 30196 53576 30248 53582
rect 30196 53518 30248 53524
rect 32864 53576 32916 53582
rect 32864 53518 32916 53524
rect 33324 53576 33376 53582
rect 33324 53518 33376 53524
rect 28632 53440 28684 53446
rect 28632 53382 28684 53388
rect 29000 53440 29052 53446
rect 29000 53382 29052 53388
rect 27528 52420 27580 52426
rect 27528 52362 27580 52368
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 29012 8090 29040 53382
rect 33704 53242 33732 53654
rect 33692 53236 33744 53242
rect 33692 53178 33744 53184
rect 34532 52426 34560 56782
rect 34624 56370 34652 57326
rect 34612 56364 34664 56370
rect 34612 56306 34664 56312
rect 34624 55350 34652 56306
rect 34612 55344 34664 55350
rect 34612 55286 34664 55292
rect 34624 54670 34652 55286
rect 34612 54664 34664 54670
rect 34612 54606 34664 54612
rect 34624 54330 34652 54606
rect 34612 54324 34664 54330
rect 34612 54266 34664 54272
rect 34624 53990 34652 54266
rect 34612 53984 34664 53990
rect 34612 53926 34664 53932
rect 34716 53242 34744 57394
rect 34796 57248 34848 57254
rect 34796 57190 34848 57196
rect 34808 56506 34836 57190
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 35072 56840 35124 56846
rect 35072 56782 35124 56788
rect 35084 56710 35112 56782
rect 35164 56772 35216 56778
rect 35164 56714 35216 56720
rect 35072 56704 35124 56710
rect 35072 56646 35124 56652
rect 35176 56506 35204 56714
rect 34796 56500 34848 56506
rect 34796 56442 34848 56448
rect 35164 56500 35216 56506
rect 35164 56442 35216 56448
rect 34808 55842 34836 56442
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34808 55814 34928 55842
rect 34796 55752 34848 55758
rect 34796 55694 34848 55700
rect 34808 54874 34836 55694
rect 34900 55146 34928 55814
rect 34980 55820 35032 55826
rect 34980 55762 35032 55768
rect 34992 55418 35020 55762
rect 35164 55616 35216 55622
rect 35164 55558 35216 55564
rect 35176 55418 35204 55558
rect 34980 55412 35032 55418
rect 34980 55354 35032 55360
rect 35164 55412 35216 55418
rect 35164 55354 35216 55360
rect 35176 55282 35204 55354
rect 35164 55276 35216 55282
rect 35164 55218 35216 55224
rect 34888 55140 34940 55146
rect 34888 55082 34940 55088
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 35360 54874 35388 59214
rect 35438 59200 35494 60000
rect 35898 59200 35954 60000
rect 36358 59200 36414 60000
rect 36818 59200 36874 60000
rect 37278 59200 37334 60000
rect 37738 59200 37794 60000
rect 38198 59200 38254 60000
rect 38658 59200 38714 60000
rect 39118 59200 39174 60000
rect 39578 59200 39634 60000
rect 40038 59200 40094 60000
rect 40498 59200 40554 60000
rect 40958 59200 41014 60000
rect 41418 59200 41474 60000
rect 41878 59200 41934 60000
rect 42338 59200 42394 60000
rect 42798 59200 42854 60000
rect 43258 59200 43314 60000
rect 43718 59200 43774 60000
rect 44178 59200 44234 60000
rect 44638 59200 44694 60000
rect 45098 59200 45154 60000
rect 45558 59200 45614 60000
rect 46018 59200 46074 60000
rect 46478 59200 46534 60000
rect 46938 59200 46994 60000
rect 47398 59200 47454 60000
rect 47858 59200 47914 60000
rect 48318 59200 48374 60000
rect 48778 59200 48834 60000
rect 49238 59200 49294 60000
rect 49698 59200 49754 60000
rect 50158 59200 50214 60000
rect 50618 59200 50674 60000
rect 51078 59200 51134 60000
rect 51538 59200 51594 60000
rect 51998 59200 52054 60000
rect 52458 59200 52514 60000
rect 52918 59200 52974 60000
rect 53378 59200 53434 60000
rect 53838 59200 53894 60000
rect 54298 59200 54354 60000
rect 54758 59200 54814 60000
rect 55218 59200 55274 60000
rect 55678 59200 55734 60000
rect 56138 59200 56194 60000
rect 35452 57338 35480 59200
rect 35624 57588 35676 57594
rect 35624 57530 35676 57536
rect 35636 57458 35664 57530
rect 35912 57458 35940 59200
rect 35624 57452 35676 57458
rect 35624 57394 35676 57400
rect 35808 57452 35860 57458
rect 35808 57394 35860 57400
rect 35900 57452 35952 57458
rect 35900 57394 35952 57400
rect 35452 57310 35664 57338
rect 35532 57248 35584 57254
rect 35532 57190 35584 57196
rect 35544 56930 35572 57190
rect 35452 56902 35572 56930
rect 35452 55418 35480 56902
rect 35532 56840 35584 56846
rect 35532 56782 35584 56788
rect 35544 56370 35572 56782
rect 35532 56364 35584 56370
rect 35532 56306 35584 56312
rect 35544 55894 35572 56306
rect 35532 55888 35584 55894
rect 35532 55830 35584 55836
rect 35440 55412 35492 55418
rect 35440 55354 35492 55360
rect 34796 54868 34848 54874
rect 34796 54810 34848 54816
rect 35348 54868 35400 54874
rect 35348 54810 35400 54816
rect 35452 54330 35480 55354
rect 35636 55350 35664 57310
rect 35716 56908 35768 56914
rect 35716 56850 35768 56856
rect 35728 56438 35756 56850
rect 35820 56522 35848 57394
rect 36084 56704 36136 56710
rect 36084 56646 36136 56652
rect 36176 56704 36228 56710
rect 36176 56646 36228 56652
rect 36096 56545 36124 56646
rect 36082 56536 36138 56545
rect 35820 56494 35940 56522
rect 35716 56432 35768 56438
rect 35716 56374 35768 56380
rect 35716 56160 35768 56166
rect 35716 56102 35768 56108
rect 35624 55344 35676 55350
rect 35624 55286 35676 55292
rect 35728 55282 35756 56102
rect 35532 55276 35584 55282
rect 35532 55218 35584 55224
rect 35716 55276 35768 55282
rect 35716 55218 35768 55224
rect 34980 54324 35032 54330
rect 34980 54266 35032 54272
rect 35440 54324 35492 54330
rect 35440 54266 35492 54272
rect 34992 54194 35020 54266
rect 34980 54188 35032 54194
rect 34980 54130 35032 54136
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 35544 53786 35572 55218
rect 35716 55140 35768 55146
rect 35716 55082 35768 55088
rect 35728 54738 35756 55082
rect 35716 54732 35768 54738
rect 35716 54674 35768 54680
rect 35728 54194 35756 54674
rect 35716 54188 35768 54194
rect 35716 54130 35768 54136
rect 35912 53786 35940 56494
rect 36082 56471 36138 56480
rect 36188 56420 36216 56646
rect 36096 56392 36216 56420
rect 36096 55758 36124 56392
rect 36084 55752 36136 55758
rect 36084 55694 36136 55700
rect 36372 54874 36400 59200
rect 36452 56840 36504 56846
rect 36452 56782 36504 56788
rect 36728 56840 36780 56846
rect 36728 56782 36780 56788
rect 36464 56506 36492 56782
rect 36544 56772 36596 56778
rect 36544 56714 36596 56720
rect 36452 56500 36504 56506
rect 36452 56442 36504 56448
rect 36556 56370 36584 56714
rect 36740 56370 36768 56782
rect 36832 56506 36860 59200
rect 37292 57458 37320 59200
rect 37188 57452 37240 57458
rect 37188 57394 37240 57400
rect 37280 57452 37332 57458
rect 37280 57394 37332 57400
rect 36820 56500 36872 56506
rect 36820 56442 36872 56448
rect 36544 56364 36596 56370
rect 36544 56306 36596 56312
rect 36728 56364 36780 56370
rect 36728 56306 36780 56312
rect 36636 56160 36688 56166
rect 36636 56102 36688 56108
rect 36648 55826 36676 56102
rect 36740 55962 36768 56306
rect 36728 55956 36780 55962
rect 36728 55898 36780 55904
rect 36636 55820 36688 55826
rect 36636 55762 36688 55768
rect 36544 55752 36596 55758
rect 36544 55694 36596 55700
rect 36556 55418 36584 55694
rect 36544 55412 36596 55418
rect 36544 55354 36596 55360
rect 36450 55312 36506 55321
rect 36450 55247 36452 55256
rect 36504 55247 36506 55256
rect 36452 55218 36504 55224
rect 36360 54868 36412 54874
rect 36360 54810 36412 54816
rect 36464 54330 36492 55218
rect 37200 54330 37228 57394
rect 37278 55720 37334 55729
rect 37278 55655 37334 55664
rect 37292 55078 37320 55655
rect 37280 55072 37332 55078
rect 37280 55014 37332 55020
rect 37292 54874 37320 55014
rect 37752 54874 37780 59200
rect 37924 56840 37976 56846
rect 37924 56782 37976 56788
rect 38108 56840 38160 56846
rect 38108 56782 38160 56788
rect 37936 55962 37964 56782
rect 37924 55956 37976 55962
rect 37924 55898 37976 55904
rect 37936 55758 37964 55898
rect 37924 55752 37976 55758
rect 37924 55694 37976 55700
rect 38120 55622 38148 56782
rect 38108 55616 38160 55622
rect 38108 55558 38160 55564
rect 37280 54868 37332 54874
rect 37280 54810 37332 54816
rect 37740 54868 37792 54874
rect 37740 54810 37792 54816
rect 36452 54324 36504 54330
rect 36452 54266 36504 54272
rect 37188 54324 37240 54330
rect 37188 54266 37240 54272
rect 34888 53780 34940 53786
rect 34888 53722 34940 53728
rect 35532 53780 35584 53786
rect 35532 53722 35584 53728
rect 35900 53780 35952 53786
rect 35900 53722 35952 53728
rect 34704 53236 34756 53242
rect 34704 53178 34756 53184
rect 34900 53174 34928 53722
rect 36464 53718 36492 54266
rect 38212 54194 38240 59200
rect 38476 57452 38528 57458
rect 38476 57394 38528 57400
rect 38292 56908 38344 56914
rect 38292 56850 38344 56856
rect 38304 56234 38332 56850
rect 38292 56228 38344 56234
rect 38292 56170 38344 56176
rect 38304 55962 38332 56170
rect 38292 55956 38344 55962
rect 38292 55898 38344 55904
rect 38384 55888 38436 55894
rect 38384 55830 38436 55836
rect 38292 55752 38344 55758
rect 38292 55694 38344 55700
rect 38304 55264 38332 55694
rect 38396 55418 38424 55830
rect 38384 55412 38436 55418
rect 38384 55354 38436 55360
rect 38384 55276 38436 55282
rect 38304 55236 38384 55264
rect 38384 55218 38436 55224
rect 38488 54874 38516 57394
rect 38672 56828 38700 59200
rect 38752 56840 38804 56846
rect 38672 56800 38752 56828
rect 38752 56782 38804 56788
rect 39026 56808 39082 56817
rect 38568 56296 38620 56302
rect 38568 56238 38620 56244
rect 38580 55894 38608 56238
rect 38568 55888 38620 55894
rect 38568 55830 38620 55836
rect 38660 55752 38712 55758
rect 38660 55694 38712 55700
rect 38672 55350 38700 55694
rect 38660 55344 38712 55350
rect 38660 55286 38712 55292
rect 38476 54868 38528 54874
rect 38476 54810 38528 54816
rect 38764 54602 38792 56782
rect 39026 56743 39082 56752
rect 39040 56438 39068 56743
rect 39132 56545 39160 59200
rect 39118 56536 39174 56545
rect 39118 56471 39174 56480
rect 39028 56432 39080 56438
rect 39028 56374 39080 56380
rect 38936 56296 38988 56302
rect 38936 56238 38988 56244
rect 38948 55894 38976 56238
rect 38936 55888 38988 55894
rect 38936 55830 38988 55836
rect 38752 54596 38804 54602
rect 38752 54538 38804 54544
rect 39040 54330 39068 56374
rect 39592 56273 39620 59200
rect 39948 57792 40000 57798
rect 39948 57734 40000 57740
rect 39960 57594 39988 57734
rect 39948 57588 40000 57594
rect 39948 57530 40000 57536
rect 39578 56264 39634 56273
rect 39578 56199 39634 56208
rect 39856 56160 39908 56166
rect 39856 56102 39908 56108
rect 39302 55992 39358 56001
rect 39302 55927 39358 55936
rect 39316 55758 39344 55927
rect 39868 55865 39896 56102
rect 39854 55856 39910 55865
rect 39854 55791 39910 55800
rect 39304 55752 39356 55758
rect 39304 55694 39356 55700
rect 39488 55752 39540 55758
rect 39488 55694 39540 55700
rect 39948 55752 40000 55758
rect 39948 55694 40000 55700
rect 39120 55684 39172 55690
rect 39120 55626 39172 55632
rect 39132 55418 39160 55626
rect 39120 55412 39172 55418
rect 39120 55354 39172 55360
rect 39316 55214 39344 55694
rect 39500 55282 39528 55694
rect 39960 55350 39988 55694
rect 39948 55344 40000 55350
rect 39948 55286 40000 55292
rect 39488 55276 39540 55282
rect 39488 55218 39540 55224
rect 39856 55276 39908 55282
rect 39856 55218 39908 55224
rect 39304 55208 39356 55214
rect 39304 55150 39356 55156
rect 39212 54664 39264 54670
rect 39316 54652 39344 55150
rect 39500 54806 39528 55218
rect 39488 54800 39540 54806
rect 39488 54742 39540 54748
rect 39868 54738 39896 55218
rect 39960 54874 39988 55286
rect 39948 54868 40000 54874
rect 39948 54810 40000 54816
rect 39856 54732 39908 54738
rect 39856 54674 39908 54680
rect 39264 54624 39344 54652
rect 39212 54606 39264 54612
rect 39028 54324 39080 54330
rect 39028 54266 39080 54272
rect 40052 54194 40080 59200
rect 40512 57474 40540 59200
rect 40512 57446 40632 57474
rect 40224 57384 40276 57390
rect 40500 57384 40552 57390
rect 40276 57344 40356 57372
rect 40224 57326 40276 57332
rect 40224 57248 40276 57254
rect 40224 57190 40276 57196
rect 40236 56914 40264 57190
rect 40328 56982 40356 57344
rect 40500 57326 40552 57332
rect 40512 57050 40540 57326
rect 40500 57044 40552 57050
rect 40500 56986 40552 56992
rect 40316 56976 40368 56982
rect 40316 56918 40368 56924
rect 40224 56908 40276 56914
rect 40224 56850 40276 56856
rect 40236 56681 40264 56850
rect 40328 56710 40356 56918
rect 40316 56704 40368 56710
rect 40222 56672 40278 56681
rect 40316 56646 40368 56652
rect 40222 56607 40278 56616
rect 40236 56370 40264 56607
rect 40224 56364 40276 56370
rect 40224 56306 40276 56312
rect 40236 55350 40264 56306
rect 40224 55344 40276 55350
rect 40224 55286 40276 55292
rect 40236 54262 40264 55286
rect 40328 55078 40356 56646
rect 40500 56296 40552 56302
rect 40500 56238 40552 56244
rect 40408 55888 40460 55894
rect 40408 55830 40460 55836
rect 40420 55690 40448 55830
rect 40408 55684 40460 55690
rect 40408 55626 40460 55632
rect 40512 55418 40540 56238
rect 40604 55826 40632 57446
rect 40684 57452 40736 57458
rect 40684 57394 40736 57400
rect 40696 56846 40724 57394
rect 40776 57044 40828 57050
rect 40776 56986 40828 56992
rect 40684 56840 40736 56846
rect 40684 56782 40736 56788
rect 40696 56302 40724 56782
rect 40684 56296 40736 56302
rect 40684 56238 40736 56244
rect 40684 56160 40736 56166
rect 40684 56102 40736 56108
rect 40592 55820 40644 55826
rect 40592 55762 40644 55768
rect 40696 55706 40724 56102
rect 40788 55894 40816 56986
rect 40868 56364 40920 56370
rect 40868 56306 40920 56312
rect 40880 55962 40908 56306
rect 40868 55956 40920 55962
rect 40868 55898 40920 55904
rect 40972 55894 41000 59200
rect 41432 57798 41460 59200
rect 41420 57792 41472 57798
rect 41420 57734 41472 57740
rect 41052 57248 41104 57254
rect 41052 57190 41104 57196
rect 41696 57248 41748 57254
rect 41696 57190 41748 57196
rect 41064 56506 41092 57190
rect 41510 56944 41566 56953
rect 41510 56879 41566 56888
rect 41604 56908 41656 56914
rect 41328 56856 41380 56862
rect 41156 56804 41328 56828
rect 41156 56800 41380 56804
rect 41052 56500 41104 56506
rect 41052 56442 41104 56448
rect 41050 56400 41106 56409
rect 41050 56335 41052 56344
rect 41104 56335 41106 56344
rect 41052 56306 41104 56312
rect 41156 56302 41184 56800
rect 41328 56798 41380 56800
rect 41524 56778 41552 56879
rect 41604 56850 41656 56856
rect 41616 56817 41644 56850
rect 41602 56808 41658 56817
rect 41512 56772 41564 56778
rect 41602 56743 41658 56752
rect 41512 56714 41564 56720
rect 41420 56704 41472 56710
rect 41418 56672 41420 56681
rect 41472 56672 41474 56681
rect 41418 56607 41474 56616
rect 41432 56302 41460 56607
rect 41616 56302 41644 56743
rect 41708 56438 41736 57190
rect 41696 56432 41748 56438
rect 41696 56374 41748 56380
rect 41144 56296 41196 56302
rect 41144 56238 41196 56244
rect 41420 56296 41472 56302
rect 41420 56238 41472 56244
rect 41604 56296 41656 56302
rect 41604 56238 41656 56244
rect 40776 55888 40828 55894
rect 40776 55830 40828 55836
rect 40960 55888 41012 55894
rect 40960 55830 41012 55836
rect 40868 55752 40920 55758
rect 40604 55690 40816 55706
rect 40868 55694 40920 55700
rect 40592 55684 40816 55690
rect 40644 55678 40816 55684
rect 40592 55626 40644 55632
rect 40788 55622 40816 55678
rect 40684 55616 40736 55622
rect 40684 55558 40736 55564
rect 40776 55616 40828 55622
rect 40776 55558 40828 55564
rect 40696 55418 40724 55558
rect 40500 55412 40552 55418
rect 40500 55354 40552 55360
rect 40684 55412 40736 55418
rect 40684 55354 40736 55360
rect 40316 55072 40368 55078
rect 40316 55014 40368 55020
rect 40328 54330 40356 55014
rect 40880 54738 40908 55694
rect 41156 55214 41184 56238
rect 41420 56160 41472 56166
rect 41420 56102 41472 56108
rect 41328 55684 41380 55690
rect 41328 55626 41380 55632
rect 41236 55412 41288 55418
rect 41340 55400 41368 55626
rect 41288 55372 41368 55400
rect 41236 55354 41288 55360
rect 41144 55208 41196 55214
rect 41144 55150 41196 55156
rect 41236 55072 41288 55078
rect 41236 55014 41288 55020
rect 40868 54732 40920 54738
rect 40868 54674 40920 54680
rect 41248 54670 41276 55014
rect 41236 54664 41288 54670
rect 41236 54606 41288 54612
rect 40316 54324 40368 54330
rect 40316 54266 40368 54272
rect 40224 54256 40276 54262
rect 40224 54198 40276 54204
rect 38200 54188 38252 54194
rect 38200 54130 38252 54136
rect 40040 54188 40092 54194
rect 40040 54130 40092 54136
rect 40052 53786 40080 54130
rect 40040 53780 40092 53786
rect 40040 53722 40092 53728
rect 36452 53712 36504 53718
rect 36452 53654 36504 53660
rect 40236 53650 40264 54198
rect 41248 54126 41276 54606
rect 41432 54330 41460 56102
rect 41696 55888 41748 55894
rect 41696 55830 41748 55836
rect 41604 55072 41656 55078
rect 41604 55014 41656 55020
rect 41420 54324 41472 54330
rect 41420 54266 41472 54272
rect 41616 54194 41644 55014
rect 41708 54874 41736 55830
rect 41892 55214 41920 59200
rect 42156 57588 42208 57594
rect 42156 57530 42208 57536
rect 42168 56846 42196 57530
rect 42156 56840 42208 56846
rect 42156 56782 42208 56788
rect 42168 56370 42196 56782
rect 42156 56364 42208 56370
rect 42156 56306 42208 56312
rect 42248 56364 42300 56370
rect 42248 56306 42300 56312
rect 42260 55894 42288 56306
rect 42248 55888 42300 55894
rect 42248 55830 42300 55836
rect 42352 55282 42380 59200
rect 42812 57458 42840 59200
rect 42800 57452 42852 57458
rect 42800 57394 42852 57400
rect 43076 57384 43128 57390
rect 43076 57326 43128 57332
rect 42432 56704 42484 56710
rect 42432 56646 42484 56652
rect 42616 56704 42668 56710
rect 42616 56646 42668 56652
rect 42444 55418 42472 56646
rect 42524 56364 42576 56370
rect 42524 56306 42576 56312
rect 42536 55962 42564 56306
rect 42524 55956 42576 55962
rect 42524 55898 42576 55904
rect 42628 55758 42656 56646
rect 43088 56370 43116 57326
rect 43168 56840 43220 56846
rect 43168 56782 43220 56788
rect 43180 56438 43208 56782
rect 43272 56506 43300 59200
rect 43352 57588 43404 57594
rect 43352 57530 43404 57536
rect 43364 57390 43392 57530
rect 43352 57384 43404 57390
rect 43352 57326 43404 57332
rect 43260 56500 43312 56506
rect 43260 56442 43312 56448
rect 43364 56438 43392 57326
rect 43732 56438 43760 59200
rect 44088 57452 44140 57458
rect 44088 57394 44140 57400
rect 43996 57316 44048 57322
rect 43996 57258 44048 57264
rect 43812 56976 43864 56982
rect 43810 56944 43812 56953
rect 43864 56944 43866 56953
rect 43810 56879 43866 56888
rect 43904 56908 43956 56914
rect 43904 56850 43956 56856
rect 43916 56817 43944 56850
rect 44008 56846 44036 57258
rect 43996 56840 44048 56846
rect 43902 56808 43958 56817
rect 43996 56782 44048 56788
rect 43902 56743 43958 56752
rect 43168 56432 43220 56438
rect 43168 56374 43220 56380
rect 43352 56432 43404 56438
rect 43352 56374 43404 56380
rect 43720 56432 43772 56438
rect 43720 56374 43772 56380
rect 43076 56364 43128 56370
rect 43076 56306 43128 56312
rect 42892 56160 42944 56166
rect 42892 56102 42944 56108
rect 42800 55888 42852 55894
rect 42800 55830 42852 55836
rect 42812 55758 42840 55830
rect 42616 55752 42668 55758
rect 42616 55694 42668 55700
rect 42800 55752 42852 55758
rect 42800 55694 42852 55700
rect 42432 55412 42484 55418
rect 42432 55354 42484 55360
rect 41972 55276 42024 55282
rect 41972 55218 42024 55224
rect 42340 55276 42392 55282
rect 42340 55218 42392 55224
rect 41880 55208 41932 55214
rect 41880 55150 41932 55156
rect 41880 55072 41932 55078
rect 41880 55014 41932 55020
rect 41696 54868 41748 54874
rect 41696 54810 41748 54816
rect 41892 54738 41920 55014
rect 41880 54732 41932 54738
rect 41880 54674 41932 54680
rect 41604 54188 41656 54194
rect 41604 54130 41656 54136
rect 41236 54120 41288 54126
rect 41236 54062 41288 54068
rect 41892 53786 41920 54674
rect 41984 54602 42012 55218
rect 41972 54596 42024 54602
rect 41972 54538 42024 54544
rect 41984 54330 42012 54538
rect 42432 54528 42484 54534
rect 42432 54470 42484 54476
rect 41972 54324 42024 54330
rect 41972 54266 42024 54272
rect 42064 54256 42116 54262
rect 42064 54198 42116 54204
rect 42076 53786 42104 54198
rect 42444 54194 42472 54470
rect 42432 54188 42484 54194
rect 42432 54130 42484 54136
rect 42248 54120 42300 54126
rect 42248 54062 42300 54068
rect 41880 53780 41932 53786
rect 41880 53722 41932 53728
rect 42064 53780 42116 53786
rect 42064 53722 42116 53728
rect 40224 53644 40276 53650
rect 40224 53586 40276 53592
rect 40776 53644 40828 53650
rect 40776 53586 40828 53592
rect 40788 53242 40816 53586
rect 42260 53514 42288 54062
rect 42248 53508 42300 53514
rect 42248 53450 42300 53456
rect 42444 53446 42472 54130
rect 42628 54126 42656 55694
rect 42708 55140 42760 55146
rect 42708 55082 42760 55088
rect 42720 54670 42748 55082
rect 42708 54664 42760 54670
rect 42708 54606 42760 54612
rect 42720 54126 42748 54606
rect 42812 54534 42840 55694
rect 42904 55622 42932 56102
rect 43088 56001 43116 56306
rect 43074 55992 43130 56001
rect 43180 55962 43208 56374
rect 44008 56370 44036 56782
rect 43536 56364 43588 56370
rect 43536 56306 43588 56312
rect 43996 56364 44048 56370
rect 43996 56306 44048 56312
rect 43074 55927 43130 55936
rect 43168 55956 43220 55962
rect 43168 55898 43220 55904
rect 43548 55826 43576 56306
rect 43536 55820 43588 55826
rect 43536 55762 43588 55768
rect 42892 55616 42944 55622
rect 42892 55558 42944 55564
rect 43548 54670 43576 55762
rect 44008 55758 44036 56306
rect 43996 55752 44048 55758
rect 43996 55694 44048 55700
rect 44100 55418 44128 57394
rect 44192 57338 44220 59200
rect 44192 57310 44312 57338
rect 44180 57248 44232 57254
rect 44180 57190 44232 57196
rect 44192 56545 44220 57190
rect 44178 56536 44234 56545
rect 44178 56471 44234 56480
rect 44284 55894 44312 57310
rect 44548 56296 44600 56302
rect 44548 56238 44600 56244
rect 44560 55962 44588 56238
rect 44652 56234 44680 59200
rect 45008 57384 45060 57390
rect 45008 57326 45060 57332
rect 44824 57248 44876 57254
rect 44824 57190 44876 57196
rect 44916 57248 44968 57254
rect 44916 57190 44968 57196
rect 44836 56273 44864 57190
rect 44822 56264 44878 56273
rect 44640 56228 44692 56234
rect 44822 56199 44878 56208
rect 44640 56170 44692 56176
rect 44548 55956 44600 55962
rect 44548 55898 44600 55904
rect 44272 55888 44324 55894
rect 44272 55830 44324 55836
rect 44560 55758 44588 55898
rect 44928 55758 44956 57190
rect 45020 55894 45048 57326
rect 45112 56302 45140 59200
rect 45192 57792 45244 57798
rect 45192 57734 45244 57740
rect 45204 56846 45232 57734
rect 45572 57526 45600 59200
rect 45560 57520 45612 57526
rect 45560 57462 45612 57468
rect 45468 57452 45520 57458
rect 45468 57394 45520 57400
rect 45480 56982 45508 57394
rect 45468 56976 45520 56982
rect 45468 56918 45520 56924
rect 45192 56840 45244 56846
rect 45192 56782 45244 56788
rect 45100 56296 45152 56302
rect 45100 56238 45152 56244
rect 45008 55888 45060 55894
rect 45008 55830 45060 55836
rect 44548 55752 44600 55758
rect 44548 55694 44600 55700
rect 44916 55752 44968 55758
rect 44916 55694 44968 55700
rect 44732 55684 44784 55690
rect 44732 55626 44784 55632
rect 44088 55412 44140 55418
rect 44088 55354 44140 55360
rect 44744 54670 44772 55626
rect 44928 54738 44956 55694
rect 45020 54874 45048 55830
rect 45204 55418 45232 56782
rect 45480 56370 45508 56918
rect 45468 56364 45520 56370
rect 45468 56306 45520 56312
rect 45468 56160 45520 56166
rect 45468 56102 45520 56108
rect 45480 55758 45508 56102
rect 45468 55752 45520 55758
rect 45468 55694 45520 55700
rect 45572 55418 45600 57462
rect 46032 56982 46060 59200
rect 46388 57248 46440 57254
rect 46388 57190 46440 57196
rect 46020 56976 46072 56982
rect 46020 56918 46072 56924
rect 46204 56840 46256 56846
rect 46204 56782 46256 56788
rect 46216 56438 46244 56782
rect 46400 56506 46428 57190
rect 46388 56500 46440 56506
rect 46388 56442 46440 56448
rect 46204 56432 46256 56438
rect 46204 56374 46256 56380
rect 46492 56370 46520 59200
rect 46952 57458 46980 59200
rect 46940 57452 46992 57458
rect 46940 57394 46992 57400
rect 46756 56840 46808 56846
rect 46756 56782 46808 56788
rect 45652 56364 45704 56370
rect 45652 56306 45704 56312
rect 46480 56364 46532 56370
rect 46480 56306 46532 56312
rect 45664 55894 45692 56306
rect 46768 55962 46796 56782
rect 46952 55962 46980 57394
rect 47412 57050 47440 59200
rect 47492 57384 47544 57390
rect 47492 57326 47544 57332
rect 47400 57044 47452 57050
rect 47400 56986 47452 56992
rect 46756 55956 46808 55962
rect 46756 55898 46808 55904
rect 46940 55956 46992 55962
rect 46940 55898 46992 55904
rect 45652 55888 45704 55894
rect 45652 55830 45704 55836
rect 45192 55412 45244 55418
rect 45192 55354 45244 55360
rect 45560 55412 45612 55418
rect 45560 55354 45612 55360
rect 45664 55350 45692 55830
rect 47504 55826 47532 57326
rect 47872 56914 47900 59200
rect 48332 57458 48360 59200
rect 48320 57452 48372 57458
rect 48320 57394 48372 57400
rect 47860 56908 47912 56914
rect 47860 56850 47912 56856
rect 48332 56506 48360 57394
rect 48792 57050 48820 59200
rect 48780 57044 48832 57050
rect 48780 56986 48832 56992
rect 49252 56982 49280 59200
rect 49712 57458 49740 59200
rect 49700 57452 49752 57458
rect 49700 57394 49752 57400
rect 49240 56976 49292 56982
rect 49240 56918 49292 56924
rect 49712 56506 49740 57394
rect 50172 57050 50200 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 50160 57044 50212 57050
rect 50160 56986 50212 56992
rect 50632 56982 50660 59200
rect 51092 57458 51120 59200
rect 51080 57452 51132 57458
rect 51080 57394 51132 57400
rect 50620 56976 50672 56982
rect 50620 56918 50672 56924
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 51092 56506 51120 57394
rect 51552 57050 51580 59200
rect 51632 57248 51684 57254
rect 51632 57190 51684 57196
rect 51540 57044 51592 57050
rect 51540 56986 51592 56992
rect 48320 56500 48372 56506
rect 48320 56442 48372 56448
rect 49700 56500 49752 56506
rect 49700 56442 49752 56448
rect 51080 56500 51132 56506
rect 51080 56442 51132 56448
rect 47492 55820 47544 55826
rect 47492 55762 47544 55768
rect 51644 55729 51672 57190
rect 52012 56982 52040 59200
rect 52472 57526 52500 59200
rect 52460 57520 52512 57526
rect 52460 57462 52512 57468
rect 52000 56976 52052 56982
rect 52000 56918 52052 56924
rect 52472 56506 52500 57462
rect 52932 57458 52960 59200
rect 52920 57452 52972 57458
rect 52920 57394 52972 57400
rect 52736 57248 52788 57254
rect 52736 57190 52788 57196
rect 52460 56500 52512 56506
rect 52460 56442 52512 56448
rect 51630 55720 51686 55729
rect 51630 55655 51686 55664
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 45652 55344 45704 55350
rect 52748 55321 52776 57190
rect 53392 57050 53420 59200
rect 53852 57458 53880 59200
rect 53840 57452 53892 57458
rect 53840 57394 53892 57400
rect 54208 57452 54260 57458
rect 54208 57394 54260 57400
rect 53380 57044 53432 57050
rect 53380 56986 53432 56992
rect 54220 56506 54248 57394
rect 54312 57050 54340 59200
rect 54772 57050 54800 59200
rect 55232 57458 55260 59200
rect 55692 57458 55720 59200
rect 55220 57452 55272 57458
rect 55220 57394 55272 57400
rect 55680 57452 55732 57458
rect 55680 57394 55732 57400
rect 55232 57050 55260 57394
rect 55404 57248 55456 57254
rect 55404 57190 55456 57196
rect 54300 57044 54352 57050
rect 54300 56986 54352 56992
rect 54760 57044 54812 57050
rect 54760 56986 54812 56992
rect 55220 57044 55272 57050
rect 55220 56986 55272 56992
rect 54208 56500 54260 56506
rect 54208 56442 54260 56448
rect 55416 55894 55444 57190
rect 56152 57050 56180 59200
rect 56140 57044 56192 57050
rect 56140 56986 56192 56992
rect 55404 55888 55456 55894
rect 55404 55830 55456 55836
rect 45652 55286 45704 55292
rect 52734 55312 52790 55321
rect 52734 55247 52790 55256
rect 45008 54868 45060 54874
rect 45008 54810 45060 54816
rect 44916 54732 44968 54738
rect 44916 54674 44968 54680
rect 43536 54664 43588 54670
rect 43536 54606 43588 54612
rect 44732 54664 44784 54670
rect 44732 54606 44784 54612
rect 42800 54528 42852 54534
rect 42800 54470 42852 54476
rect 44180 54528 44232 54534
rect 44180 54470 44232 54476
rect 44192 54194 44220 54470
rect 44744 54262 44772 54606
rect 44732 54256 44784 54262
rect 44732 54198 44784 54204
rect 44180 54188 44232 54194
rect 44180 54130 44232 54136
rect 44928 54126 44956 54674
rect 45020 54194 45048 54810
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 45008 54188 45060 54194
rect 45008 54130 45060 54136
rect 42616 54120 42668 54126
rect 42616 54062 42668 54068
rect 42708 54120 42760 54126
rect 42708 54062 42760 54068
rect 44916 54120 44968 54126
rect 44916 54062 44968 54068
rect 42432 53440 42484 53446
rect 42432 53382 42484 53388
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 40776 53236 40828 53242
rect 40776 53178 40828 53184
rect 34888 53168 34940 53174
rect 34888 53110 34940 53116
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34520 52420 34572 52426
rect 34520 52362 34572 52368
rect 34532 52086 34560 52362
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 34520 52080 34572 52086
rect 34520 52022 34572 52028
rect 34060 51944 34112 51950
rect 34060 51886 34112 51892
rect 35808 51944 35860 51950
rect 35808 51886 35860 51892
rect 34072 51610 34100 51886
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34060 51604 34112 51610
rect 34060 51546 34112 51552
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 29000 8084 29052 8090
rect 29000 8026 29052 8032
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 29012 7426 29040 8026
rect 29564 7954 29592 8434
rect 30196 8356 30248 8362
rect 30196 8298 30248 8304
rect 29552 7948 29604 7954
rect 29552 7890 29604 7896
rect 29460 7880 29512 7886
rect 29460 7822 29512 7828
rect 29012 7410 29132 7426
rect 26976 7404 27028 7410
rect 26976 7346 27028 7352
rect 29012 7404 29144 7410
rect 29012 7398 29092 7404
rect 26884 7200 26936 7206
rect 26884 7142 26936 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 26424 6656 26476 6662
rect 26424 6598 26476 6604
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 26436 6322 26464 6598
rect 26424 6316 26476 6322
rect 26424 6258 26476 6264
rect 25320 6112 25372 6118
rect 25320 6054 25372 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 25332 5234 25360 6054
rect 26436 5846 26464 6258
rect 26424 5840 26476 5846
rect 26424 5782 26476 5788
rect 26896 5778 26924 7142
rect 26988 6798 27016 7346
rect 27712 7336 27764 7342
rect 27712 7278 27764 7284
rect 27896 7336 27948 7342
rect 27896 7278 27948 7284
rect 26976 6792 27028 6798
rect 26976 6734 27028 6740
rect 27620 6792 27672 6798
rect 27620 6734 27672 6740
rect 26988 6254 27016 6734
rect 27632 6322 27660 6734
rect 27620 6316 27672 6322
rect 27620 6258 27672 6264
rect 26976 6248 27028 6254
rect 26976 6190 27028 6196
rect 27436 6248 27488 6254
rect 27436 6190 27488 6196
rect 26884 5772 26936 5778
rect 26884 5714 26936 5720
rect 25504 5568 25556 5574
rect 25504 5510 25556 5516
rect 25516 5302 25544 5510
rect 25504 5296 25556 5302
rect 25504 5238 25556 5244
rect 27448 5234 27476 6190
rect 27724 6186 27752 7278
rect 27804 6656 27856 6662
rect 27804 6598 27856 6604
rect 27816 6390 27844 6598
rect 27804 6384 27856 6390
rect 27804 6326 27856 6332
rect 27712 6180 27764 6186
rect 27712 6122 27764 6128
rect 27528 5772 27580 5778
rect 27528 5714 27580 5720
rect 25320 5228 25372 5234
rect 25320 5170 25372 5176
rect 27436 5228 27488 5234
rect 27436 5170 27488 5176
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 26240 5160 26292 5166
rect 26240 5102 26292 5108
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 7668 800 7696 2790
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8220 800 8248 2382
rect 8588 800 8616 2790
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 8956 800 8984 2382
rect 9324 800 9352 3470
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9692 800 9720 2518
rect 9968 800 9996 2790
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10244 800 10272 2382
rect 10520 800 10548 2790
rect 10796 800 10824 3470
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 11072 800 11100 2790
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 11348 800 11376 2518
rect 11624 800 11652 2790
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11900 800 11928 2382
rect 12176 800 12204 2790
rect 12452 800 12480 3470
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 12728 800 12756 2450
rect 13004 800 13032 2790
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13280 800 13308 2382
rect 13556 800 13584 3470
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 13832 800 13860 2790
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14108 800 14136 2382
rect 14384 800 14412 2790
rect 14660 800 14688 3470
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 14936 800 14964 2518
rect 15212 800 15240 2790
rect 15488 800 15516 3470
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 15752 2372 15804 2378
rect 15752 2314 15804 2320
rect 15764 800 15792 2314
rect 16040 800 16068 2790
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16316 800 16344 2382
rect 16592 800 16620 3470
rect 16856 2984 16908 2990
rect 16856 2926 16908 2932
rect 16868 800 16896 2926
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 17144 800 17172 2790
rect 17328 800 17356 3470
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 17604 800 17632 2450
rect 17880 800 17908 2790
rect 18156 800 18184 3470
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 18432 800 18460 2518
rect 18708 800 18736 2790
rect 18984 800 19012 3470
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 19260 800 19288 2450
rect 19444 1442 19472 2790
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 1986 20024 3878
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20076 2576 20128 2582
rect 20076 2518 20128 2524
rect 19812 1958 20024 1986
rect 19444 1414 19564 1442
rect 19536 800 19564 1414
rect 19812 800 19840 1958
rect 20088 800 20116 2518
rect 20364 800 20392 3470
rect 20640 800 20668 3878
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20916 800 20944 3470
rect 21180 2984 21232 2990
rect 21180 2926 21232 2932
rect 21192 800 21220 2926
rect 21468 800 21496 4558
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 21732 2916 21784 2922
rect 21732 2858 21784 2864
rect 21744 800 21772 2858
rect 22020 800 22048 3878
rect 22284 3664 22336 3670
rect 22284 3606 22336 3612
rect 22192 3528 22244 3534
rect 22192 3470 22244 3476
rect 22204 3058 22232 3470
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 22296 800 22324 3606
rect 22572 800 22600 4558
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 22848 3058 22876 3674
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 22848 800 22876 2450
rect 23124 800 23152 4966
rect 23940 4752 23992 4758
rect 23940 4694 23992 4700
rect 23664 4004 23716 4010
rect 23664 3946 23716 3952
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23400 800 23428 2926
rect 23584 2650 23612 3470
rect 23572 2644 23624 2650
rect 23572 2586 23624 2592
rect 23676 800 23704 3946
rect 23756 2372 23808 2378
rect 23756 2314 23808 2320
rect 23768 1426 23796 2314
rect 23756 1420 23808 1426
rect 23756 1362 23808 1368
rect 23952 800 23980 4694
rect 24124 4616 24176 4622
rect 24124 4558 24176 4564
rect 24136 4146 24164 4558
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 24136 3670 24164 4082
rect 24492 3936 24544 3942
rect 24492 3878 24544 3884
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 24504 3670 24532 3878
rect 24124 3664 24176 3670
rect 24124 3606 24176 3612
rect 24492 3664 24544 3670
rect 24492 3606 24544 3612
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 24216 3052 24268 3058
rect 24216 2994 24268 3000
rect 24032 2916 24084 2922
rect 24032 2858 24084 2864
rect 24044 2378 24072 2858
rect 24228 2446 24256 2994
rect 24124 2440 24176 2446
rect 24124 2382 24176 2388
rect 24216 2440 24268 2446
rect 24216 2382 24268 2388
rect 24032 2372 24084 2378
rect 24032 2314 24084 2320
rect 24136 2106 24164 2382
rect 24124 2100 24176 2106
rect 24124 2042 24176 2048
rect 24320 1170 24348 3334
rect 24688 3194 24716 3878
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24676 2984 24728 2990
rect 24674 2952 24676 2961
rect 24728 2952 24730 2961
rect 24674 2887 24730 2896
rect 24492 1420 24544 1426
rect 24492 1362 24544 1368
rect 24228 1142 24348 1170
rect 24228 800 24256 1142
rect 24504 800 24532 1362
rect 24780 800 24808 5102
rect 25872 5024 25924 5030
rect 25872 4966 25924 4972
rect 25884 4690 25912 4966
rect 25872 4684 25924 4690
rect 25872 4626 25924 4632
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 26148 4140 26200 4146
rect 26148 4082 26200 4088
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 25424 3670 25452 3878
rect 25320 3664 25372 3670
rect 25320 3606 25372 3612
rect 25412 3664 25464 3670
rect 25412 3606 25464 3612
rect 25044 2576 25096 2582
rect 25044 2518 25096 2524
rect 25056 800 25084 2518
rect 25332 800 25360 3606
rect 25516 3058 25544 4082
rect 25872 4072 25924 4078
rect 25872 4014 25924 4020
rect 25884 3534 25912 4014
rect 26160 3942 26188 4082
rect 26056 3936 26108 3942
rect 26056 3878 26108 3884
rect 26148 3936 26200 3942
rect 26148 3878 26200 3884
rect 25872 3528 25924 3534
rect 25872 3470 25924 3476
rect 26068 3398 26096 3878
rect 26056 3392 26108 3398
rect 26056 3334 26108 3340
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 25596 2984 25648 2990
rect 25596 2926 25648 2932
rect 25504 2848 25556 2854
rect 25504 2790 25556 2796
rect 25516 1442 25544 2790
rect 25608 2650 25636 2926
rect 26252 2802 26280 5102
rect 26332 5092 26384 5098
rect 26332 5034 26384 5040
rect 26344 3942 26372 5034
rect 27252 4752 27304 4758
rect 27252 4694 27304 4700
rect 26424 4684 26476 4690
rect 26424 4626 26476 4632
rect 26332 3936 26384 3942
rect 26332 3878 26384 3884
rect 26160 2774 26280 2802
rect 25596 2644 25648 2650
rect 25596 2586 25648 2592
rect 25872 2100 25924 2106
rect 25872 2042 25924 2048
rect 25516 1414 25636 1442
rect 25608 800 25636 1414
rect 25884 800 25912 2042
rect 26160 800 26188 2774
rect 26436 800 26464 4626
rect 26608 4072 26660 4078
rect 26608 4014 26660 4020
rect 26516 3936 26568 3942
rect 26516 3878 26568 3884
rect 26528 3398 26556 3878
rect 26620 3738 26648 4014
rect 26608 3732 26660 3738
rect 26608 3674 26660 3680
rect 27264 3534 27292 4694
rect 27448 4282 27476 5170
rect 27436 4276 27488 4282
rect 27436 4218 27488 4224
rect 27252 3528 27304 3534
rect 27252 3470 27304 3476
rect 26700 3460 26752 3466
rect 26700 3402 26752 3408
rect 26516 3392 26568 3398
rect 26516 3334 26568 3340
rect 26712 800 26740 3402
rect 26976 3392 27028 3398
rect 26976 3334 27028 3340
rect 26988 800 27016 3334
rect 27252 2372 27304 2378
rect 27252 2314 27304 2320
rect 27264 800 27292 2314
rect 27540 800 27568 5714
rect 27908 5370 27936 7278
rect 29012 6914 29040 7398
rect 29092 7346 29144 7352
rect 29184 7336 29236 7342
rect 29184 7278 29236 7284
rect 29012 6886 29132 6914
rect 29104 6458 29132 6886
rect 29092 6452 29144 6458
rect 29092 6394 29144 6400
rect 29104 6322 29132 6394
rect 29092 6316 29144 6322
rect 29092 6258 29144 6264
rect 28080 6248 28132 6254
rect 28080 6190 28132 6196
rect 27896 5364 27948 5370
rect 27896 5306 27948 5312
rect 27896 4820 27948 4826
rect 27896 4762 27948 4768
rect 27804 3460 27856 3466
rect 27804 3402 27856 3408
rect 27620 3052 27672 3058
rect 27620 2994 27672 3000
rect 27632 2514 27660 2994
rect 27620 2508 27672 2514
rect 27620 2450 27672 2456
rect 27816 800 27844 3402
rect 27908 3058 27936 4762
rect 27896 3052 27948 3058
rect 27896 2994 27948 3000
rect 28092 800 28120 6190
rect 28908 5704 28960 5710
rect 28908 5646 28960 5652
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 28920 5234 28948 5646
rect 28908 5228 28960 5234
rect 28908 5170 28960 5176
rect 29012 5098 29040 5646
rect 29000 5092 29052 5098
rect 29000 5034 29052 5040
rect 29012 4622 29040 5034
rect 28540 4616 28592 4622
rect 28540 4558 28592 4564
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 28552 4146 28580 4558
rect 28540 4140 28592 4146
rect 28540 4082 28592 4088
rect 28908 4004 28960 4010
rect 28908 3946 28960 3952
rect 28356 3664 28408 3670
rect 28356 3606 28408 3612
rect 28368 800 28396 3606
rect 28632 2984 28684 2990
rect 28632 2926 28684 2932
rect 28644 800 28672 2926
rect 28920 800 28948 3946
rect 29012 3602 29040 4558
rect 29000 3596 29052 3602
rect 29000 3538 29052 3544
rect 29196 3466 29224 7278
rect 29472 6866 29500 7822
rect 29564 7342 29592 7890
rect 30012 7880 30064 7886
rect 30012 7822 30064 7828
rect 29552 7336 29604 7342
rect 29552 7278 29604 7284
rect 29460 6860 29512 6866
rect 29460 6802 29512 6808
rect 29460 6724 29512 6730
rect 29460 6666 29512 6672
rect 29472 5914 29500 6666
rect 29460 5908 29512 5914
rect 29460 5850 29512 5856
rect 29564 5710 29592 7278
rect 30024 5778 30052 7822
rect 30208 5778 30236 8298
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 31208 7744 31260 7750
rect 31208 7686 31260 7692
rect 30564 6996 30616 7002
rect 30564 6938 30616 6944
rect 30288 6860 30340 6866
rect 30288 6802 30340 6808
rect 30012 5772 30064 5778
rect 30012 5714 30064 5720
rect 30196 5772 30248 5778
rect 30196 5714 30248 5720
rect 29552 5704 29604 5710
rect 29552 5646 29604 5652
rect 29736 4072 29788 4078
rect 29736 4014 29788 4020
rect 29184 3460 29236 3466
rect 29184 3402 29236 3408
rect 29184 2848 29236 2854
rect 29184 2790 29236 2796
rect 29196 800 29224 2790
rect 29460 2508 29512 2514
rect 29460 2450 29512 2456
rect 29472 800 29500 2450
rect 29748 800 29776 4014
rect 30012 2848 30064 2854
rect 30012 2790 30064 2796
rect 30024 800 30052 2790
rect 30300 800 30328 6802
rect 30576 6390 30604 6938
rect 31220 6866 31248 7686
rect 31576 7404 31628 7410
rect 31576 7346 31628 7352
rect 31300 7200 31352 7206
rect 31300 7142 31352 7148
rect 31208 6860 31260 6866
rect 31208 6802 31260 6808
rect 31312 6730 31340 7142
rect 31588 7002 31616 7346
rect 33784 7200 33836 7206
rect 33784 7142 33836 7148
rect 31576 6996 31628 7002
rect 31576 6938 31628 6944
rect 31588 6866 31616 6938
rect 31484 6860 31536 6866
rect 31484 6802 31536 6808
rect 31576 6860 31628 6866
rect 31576 6802 31628 6808
rect 31300 6724 31352 6730
rect 31300 6666 31352 6672
rect 30564 6384 30616 6390
rect 30564 6326 30616 6332
rect 30576 5930 30604 6326
rect 30484 5902 30696 5930
rect 30380 5160 30432 5166
rect 30380 5102 30432 5108
rect 30392 2854 30420 5102
rect 30484 4010 30512 5902
rect 30668 5778 30696 5902
rect 30564 5772 30616 5778
rect 30564 5714 30616 5720
rect 30656 5772 30708 5778
rect 30656 5714 30708 5720
rect 30472 4004 30524 4010
rect 30472 3946 30524 3952
rect 30484 3058 30512 3946
rect 30472 3052 30524 3058
rect 30472 2994 30524 3000
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30576 800 30604 5714
rect 30840 5296 30892 5302
rect 30840 5238 30892 5244
rect 30748 4684 30800 4690
rect 30748 4626 30800 4632
rect 30656 3460 30708 3466
rect 30656 3402 30708 3408
rect 30668 3194 30696 3402
rect 30656 3188 30708 3194
rect 30656 3130 30708 3136
rect 30760 2258 30788 4626
rect 30852 3738 30880 5238
rect 31300 5160 31352 5166
rect 31300 5102 31352 5108
rect 31312 4146 31340 5102
rect 31300 4140 31352 4146
rect 31300 4082 31352 4088
rect 31496 4026 31524 6802
rect 32588 6248 32640 6254
rect 32588 6190 32640 6196
rect 33048 6248 33100 6254
rect 33048 6190 33100 6196
rect 32496 6180 32548 6186
rect 32496 6122 32548 6128
rect 32508 5914 32536 6122
rect 32496 5908 32548 5914
rect 32496 5850 32548 5856
rect 31760 5160 31812 5166
rect 31760 5102 31812 5108
rect 31496 3998 31708 4026
rect 31484 3936 31536 3942
rect 31484 3878 31536 3884
rect 30840 3732 30892 3738
rect 30840 3674 30892 3680
rect 31496 3602 31524 3878
rect 31484 3596 31536 3602
rect 31484 3538 31536 3544
rect 31392 3052 31444 3058
rect 31392 2994 31444 3000
rect 31116 2508 31168 2514
rect 31116 2450 31168 2456
rect 30760 2230 30880 2258
rect 30852 800 30880 2230
rect 31128 800 31156 2450
rect 31404 800 31432 2994
rect 31680 800 31708 3998
rect 31772 3058 31800 5102
rect 31944 3596 31996 3602
rect 31944 3538 31996 3544
rect 31760 3052 31812 3058
rect 31760 2994 31812 3000
rect 31758 2952 31814 2961
rect 31758 2887 31814 2896
rect 31772 2514 31800 2887
rect 31760 2508 31812 2514
rect 31760 2450 31812 2456
rect 31956 800 31984 3538
rect 32600 3210 32628 6190
rect 33060 5914 33088 6190
rect 33048 5908 33100 5914
rect 33048 5850 33100 5856
rect 33796 5302 33824 7142
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35820 6914 35848 51886
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 34716 6886 35848 6914
rect 34428 6656 34480 6662
rect 34428 6598 34480 6604
rect 34244 6112 34296 6118
rect 34244 6054 34296 6060
rect 33876 5840 33928 5846
rect 33876 5782 33928 5788
rect 33784 5296 33836 5302
rect 33784 5238 33836 5244
rect 33600 5160 33652 5166
rect 33600 5102 33652 5108
rect 33612 4826 33640 5102
rect 33600 4820 33652 4826
rect 33600 4762 33652 4768
rect 33048 4072 33100 4078
rect 33048 4014 33100 4020
rect 32508 3182 32628 3210
rect 32220 2984 32272 2990
rect 32220 2926 32272 2932
rect 32232 800 32260 2926
rect 32508 800 32536 3182
rect 32772 2848 32824 2854
rect 32772 2790 32824 2796
rect 32784 800 32812 2790
rect 33060 800 33088 4014
rect 33416 3936 33468 3942
rect 33416 3878 33468 3884
rect 33232 3392 33284 3398
rect 33232 3334 33284 3340
rect 33244 3126 33272 3334
rect 33232 3120 33284 3126
rect 33232 3062 33284 3068
rect 33428 3058 33456 3878
rect 33416 3052 33468 3058
rect 33416 2994 33468 3000
rect 33324 2916 33376 2922
rect 33324 2858 33376 2864
rect 33336 800 33364 2858
rect 33600 2372 33652 2378
rect 33600 2314 33652 2320
rect 33612 800 33640 2314
rect 33888 800 33916 5782
rect 34256 5778 34284 6054
rect 34440 5778 34468 6598
rect 34244 5772 34296 5778
rect 34244 5714 34296 5720
rect 34428 5772 34480 5778
rect 34428 5714 34480 5720
rect 34060 5160 34112 5166
rect 34060 5102 34112 5108
rect 34072 2854 34100 5102
rect 34520 4616 34572 4622
rect 34520 4558 34572 4564
rect 34152 4548 34204 4554
rect 34152 4490 34204 4496
rect 34060 2848 34112 2854
rect 34060 2790 34112 2796
rect 34164 800 34192 4490
rect 34532 4146 34560 4558
rect 34520 4140 34572 4146
rect 34520 4082 34572 4088
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 34440 800 34468 3538
rect 34716 800 34744 6886
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 36084 5024 36136 5030
rect 36084 4966 36136 4972
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 36096 4690 36124 4966
rect 36084 4684 36136 4690
rect 36084 4626 36136 4632
rect 36728 4616 36780 4622
rect 36728 4558 36780 4564
rect 36740 4146 36768 4558
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 36728 4140 36780 4146
rect 36728 4082 36780 4088
rect 35716 3936 35768 3942
rect 35716 3878 35768 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35728 3058 35756 3878
rect 36084 3732 36136 3738
rect 36084 3674 36136 3680
rect 35716 3052 35768 3058
rect 35716 2994 35768 3000
rect 35348 2984 35400 2990
rect 35348 2926 35400 2932
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34980 2576 35032 2582
rect 34980 2518 35032 2524
rect 34992 800 35020 2518
rect 35360 1578 35388 2926
rect 35808 2916 35860 2922
rect 35808 2858 35860 2864
rect 35530 2816 35586 2825
rect 35530 2751 35586 2760
rect 35268 1550 35388 1578
rect 35268 800 35296 1550
rect 35544 800 35572 2751
rect 35820 800 35848 2858
rect 36096 800 36124 3674
rect 36544 3664 36596 3670
rect 36544 3606 36596 3612
rect 36176 2848 36228 2854
rect 36176 2790 36228 2796
rect 36188 2514 36216 2790
rect 36176 2508 36228 2514
rect 36176 2450 36228 2456
rect 36556 2446 36584 3606
rect 36740 3534 36768 4082
rect 37188 4004 37240 4010
rect 37188 3946 37240 3952
rect 36728 3528 36780 3534
rect 36728 3470 36780 3476
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 36740 3058 36768 3470
rect 36728 3052 36780 3058
rect 36728 2994 36780 3000
rect 36740 2446 36768 2994
rect 36544 2440 36596 2446
rect 36544 2382 36596 2388
rect 36728 2440 36780 2446
rect 36728 2382 36780 2388
rect 36360 2304 36412 2310
rect 36360 2246 36412 2252
rect 36372 800 36400 2246
rect 36832 1850 36860 3470
rect 36912 2848 36964 2854
rect 36912 2790 36964 2796
rect 36648 1822 36860 1850
rect 36648 800 36676 1822
rect 36924 800 36952 2790
rect 37200 800 37228 3946
rect 37280 3936 37332 3942
rect 37280 3878 37332 3884
rect 38568 3936 38620 3942
rect 38568 3878 38620 3884
rect 37292 3602 37320 3878
rect 37280 3596 37332 3602
rect 37280 3538 37332 3544
rect 37556 3596 37608 3602
rect 37556 3538 37608 3544
rect 37464 3460 37516 3466
rect 37464 3402 37516 3408
rect 37476 2650 37504 3402
rect 37464 2644 37516 2650
rect 37464 2586 37516 2592
rect 37568 1850 37596 3538
rect 38016 3052 38068 3058
rect 38016 2994 38068 3000
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 37476 1822 37596 1850
rect 37476 800 37504 1822
rect 37752 800 37780 2314
rect 38028 800 38056 2994
rect 38292 2576 38344 2582
rect 38292 2518 38344 2524
rect 38304 800 38332 2518
rect 38580 800 38608 3878
rect 39948 3664 40000 3670
rect 39948 3606 40000 3612
rect 39396 3528 39448 3534
rect 39396 3470 39448 3476
rect 38844 2916 38896 2922
rect 38844 2858 38896 2864
rect 38658 2816 38714 2825
rect 38658 2751 38714 2760
rect 38672 2650 38700 2751
rect 38660 2644 38712 2650
rect 38660 2586 38712 2592
rect 38856 800 38884 2858
rect 39120 2508 39172 2514
rect 39120 2450 39172 2456
rect 39132 800 39160 2450
rect 39408 800 39436 3470
rect 39672 2984 39724 2990
rect 39672 2926 39724 2932
rect 39684 800 39712 2926
rect 39960 800 39988 3606
rect 40776 3596 40828 3602
rect 40776 3538 40828 3544
rect 40224 3052 40276 3058
rect 40224 2994 40276 3000
rect 40236 800 40264 2994
rect 40500 2372 40552 2378
rect 40500 2314 40552 2320
rect 40512 800 40540 2314
rect 40788 800 40816 3538
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 42432 3528 42484 3534
rect 42432 3470 42484 3476
rect 43260 3528 43312 3534
rect 43260 3470 43312 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 46020 3528 46072 3534
rect 46020 3470 46072 3476
rect 46572 3528 46624 3534
rect 46572 3470 46624 3476
rect 48228 3528 48280 3534
rect 48228 3470 48280 3476
rect 49332 3528 49384 3534
rect 49332 3470 49384 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 52092 3528 52144 3534
rect 52092 3470 52144 3476
rect 41052 2916 41104 2922
rect 41052 2858 41104 2864
rect 41064 800 41092 2858
rect 41340 800 41368 3470
rect 41880 2848 41932 2854
rect 41880 2790 41932 2796
rect 41604 2576 41656 2582
rect 41604 2518 41656 2524
rect 41616 800 41644 2518
rect 41892 800 41920 2790
rect 42156 2508 42208 2514
rect 42156 2450 42208 2456
rect 42168 800 42196 2450
rect 42444 800 42472 3470
rect 42984 2916 43036 2922
rect 42984 2858 43036 2864
rect 42708 2440 42760 2446
rect 42708 2382 42760 2388
rect 42720 800 42748 2382
rect 42996 800 43024 2858
rect 43272 800 43300 3470
rect 43536 2848 43588 2854
rect 43536 2790 43588 2796
rect 43548 800 43576 2790
rect 43812 2372 43864 2378
rect 43812 2314 43864 2320
rect 43824 800 43852 2314
rect 44100 800 44128 3470
rect 45468 2984 45520 2990
rect 45468 2926 45520 2932
rect 44364 2916 44416 2922
rect 44364 2858 44416 2864
rect 44376 800 44404 2858
rect 44916 2848 44968 2854
rect 44916 2790 44968 2796
rect 44640 2508 44692 2514
rect 44640 2450 44692 2456
rect 44652 800 44680 2450
rect 44928 800 44956 2790
rect 45192 2576 45244 2582
rect 45192 2518 45244 2524
rect 45204 800 45232 2518
rect 45480 800 45508 2926
rect 45744 2440 45796 2446
rect 45744 2382 45796 2388
rect 45756 800 45784 2382
rect 46032 800 46060 3470
rect 46296 2848 46348 2854
rect 46296 2790 46348 2796
rect 46308 800 46336 2790
rect 46584 800 46612 3470
rect 46848 2984 46900 2990
rect 46848 2926 46900 2932
rect 46860 800 46888 2926
rect 47676 2916 47728 2922
rect 47676 2858 47728 2864
rect 47124 2508 47176 2514
rect 47124 2450 47176 2456
rect 47136 800 47164 2450
rect 47400 2372 47452 2378
rect 47400 2314 47452 2320
rect 47412 800 47440 2314
rect 47688 800 47716 2858
rect 47952 2644 48004 2650
rect 47952 2586 48004 2592
rect 47964 800 47992 2586
rect 48240 800 48268 3470
rect 49056 2916 49108 2922
rect 49056 2858 49108 2864
rect 48504 2848 48556 2854
rect 48504 2790 48556 2796
rect 48516 800 48544 2790
rect 48780 2576 48832 2582
rect 48780 2518 48832 2524
rect 48792 800 48820 2518
rect 49068 800 49096 2858
rect 49344 800 49372 3470
rect 49608 2848 49660 2854
rect 49608 2790 49660 2796
rect 49620 800 49648 2790
rect 49884 2508 49936 2514
rect 49884 2450 49936 2456
rect 49896 800 49924 2450
rect 50172 800 50200 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50988 2916 51040 2922
rect 50988 2858 51040 2864
rect 50620 2848 50672 2854
rect 50620 2790 50672 2796
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50632 1442 50660 2790
rect 50712 2576 50764 2582
rect 50712 2518 50764 2524
rect 50448 1414 50660 1442
rect 50448 800 50476 1414
rect 50724 800 50752 2518
rect 51000 800 51028 2858
rect 51540 2848 51592 2854
rect 51540 2790 51592 2796
rect 51264 2372 51316 2378
rect 51264 2314 51316 2320
rect 51276 800 51304 2314
rect 51552 800 51580 2790
rect 51816 2508 51868 2514
rect 51816 2450 51868 2456
rect 51828 800 51856 2450
rect 52104 800 52132 3470
rect 52368 2916 52420 2922
rect 52368 2858 52420 2864
rect 52380 800 52408 2858
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
<< via2 >>
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 21454 57432 21510 57488
rect 22282 56616 22338 56672
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 23294 56480 23350 56536
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 23938 57432 23994 57488
rect 25502 56364 25558 56400
rect 25502 56344 25504 56364
rect 25504 56344 25556 56364
rect 25556 56344 25558 56364
rect 26238 56616 26294 56672
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 26974 55800 27030 55856
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 29274 56788 29276 56808
rect 29276 56788 29328 56808
rect 29328 56788 29330 56808
rect 29274 56752 29330 56788
rect 29274 56480 29330 56536
rect 30654 56752 30710 56808
rect 29274 55564 29276 55584
rect 29276 55564 29328 55584
rect 29328 55564 29330 55584
rect 29274 55528 29330 55564
rect 32862 55528 32918 55584
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 36082 56480 36138 56536
rect 36450 55276 36506 55312
rect 36450 55256 36452 55276
rect 36452 55256 36504 55276
rect 36504 55256 36506 55276
rect 37278 55664 37334 55720
rect 39026 56752 39082 56808
rect 39118 56480 39174 56536
rect 39578 56208 39634 56264
rect 39302 55936 39358 55992
rect 39854 55800 39910 55856
rect 40222 56616 40278 56672
rect 41510 56888 41566 56944
rect 41050 56364 41106 56400
rect 41050 56344 41052 56364
rect 41052 56344 41104 56364
rect 41104 56344 41106 56364
rect 41602 56752 41658 56808
rect 41418 56652 41420 56672
rect 41420 56652 41472 56672
rect 41472 56652 41474 56672
rect 41418 56616 41474 56652
rect 43810 56924 43812 56944
rect 43812 56924 43864 56944
rect 43864 56924 43866 56944
rect 43810 56888 43866 56924
rect 43902 56752 43958 56808
rect 43074 55936 43130 55992
rect 44178 56480 44234 56536
rect 44822 56208 44878 56264
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 51630 55664 51686 55720
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 52734 55256 52790 55312
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 24674 2932 24676 2952
rect 24676 2932 24728 2952
rect 24728 2932 24730 2952
rect 24674 2896 24730 2932
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 31758 2896 31814 2952
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35530 2760 35586 2816
rect 38658 2760 38714 2816
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
<< metal3 >>
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 21449 57490 21515 57493
rect 23933 57490 23999 57493
rect 21449 57488 23999 57490
rect 21449 57432 21454 57488
rect 21510 57432 23938 57488
rect 23994 57432 23999 57488
rect 21449 57430 23999 57432
rect 21449 57427 21515 57430
rect 23933 57427 23999 57430
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 41505 56946 41571 56949
rect 43805 56946 43871 56949
rect 41505 56944 43871 56946
rect 41505 56888 41510 56944
rect 41566 56888 43810 56944
rect 43866 56888 43871 56944
rect 41505 56886 43871 56888
rect 41505 56883 41571 56886
rect 43805 56883 43871 56886
rect 29269 56810 29335 56813
rect 30649 56810 30715 56813
rect 29269 56808 30715 56810
rect 29269 56752 29274 56808
rect 29330 56752 30654 56808
rect 30710 56752 30715 56808
rect 29269 56750 30715 56752
rect 29269 56747 29335 56750
rect 30649 56747 30715 56750
rect 39021 56810 39087 56813
rect 41597 56810 41663 56813
rect 43897 56810 43963 56813
rect 39021 56808 43963 56810
rect 39021 56752 39026 56808
rect 39082 56752 41602 56808
rect 41658 56752 43902 56808
rect 43958 56752 43963 56808
rect 39021 56750 43963 56752
rect 39021 56747 39087 56750
rect 41597 56747 41663 56750
rect 43897 56747 43963 56750
rect 22277 56674 22343 56677
rect 26233 56674 26299 56677
rect 22277 56672 26299 56674
rect 22277 56616 22282 56672
rect 22338 56616 26238 56672
rect 26294 56616 26299 56672
rect 22277 56614 26299 56616
rect 22277 56611 22343 56614
rect 26233 56611 26299 56614
rect 40217 56674 40283 56677
rect 41413 56674 41479 56677
rect 40217 56672 41479 56674
rect 40217 56616 40222 56672
rect 40278 56616 41418 56672
rect 41474 56616 41479 56672
rect 40217 56614 41479 56616
rect 40217 56611 40283 56614
rect 41413 56611 41479 56614
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 23289 56538 23355 56541
rect 29269 56538 29335 56541
rect 36077 56538 36143 56541
rect 23289 56536 36143 56538
rect 23289 56480 23294 56536
rect 23350 56480 29274 56536
rect 29330 56480 36082 56536
rect 36138 56480 36143 56536
rect 23289 56478 36143 56480
rect 23289 56475 23355 56478
rect 29269 56475 29335 56478
rect 36077 56475 36143 56478
rect 39113 56538 39179 56541
rect 44173 56538 44239 56541
rect 39113 56536 44239 56538
rect 39113 56480 39118 56536
rect 39174 56480 44178 56536
rect 44234 56480 44239 56536
rect 39113 56478 44239 56480
rect 39113 56475 39179 56478
rect 44173 56475 44239 56478
rect 25497 56402 25563 56405
rect 41045 56402 41111 56405
rect 25497 56400 41111 56402
rect 25497 56344 25502 56400
rect 25558 56344 41050 56400
rect 41106 56344 41111 56400
rect 25497 56342 41111 56344
rect 25497 56339 25563 56342
rect 41045 56339 41111 56342
rect 39573 56266 39639 56269
rect 44817 56266 44883 56269
rect 39573 56264 44883 56266
rect 39573 56208 39578 56264
rect 39634 56208 44822 56264
rect 44878 56208 44883 56264
rect 39573 56206 44883 56208
rect 39573 56203 39639 56206
rect 44817 56203 44883 56206
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 39297 55994 39363 55997
rect 43069 55994 43135 55997
rect 39297 55992 43135 55994
rect 39297 55936 39302 55992
rect 39358 55936 43074 55992
rect 43130 55936 43135 55992
rect 39297 55934 43135 55936
rect 39297 55931 39363 55934
rect 43069 55931 43135 55934
rect 26969 55858 27035 55861
rect 39849 55858 39915 55861
rect 26969 55856 39915 55858
rect 26969 55800 26974 55856
rect 27030 55800 39854 55856
rect 39910 55800 39915 55856
rect 26969 55798 39915 55800
rect 26969 55795 27035 55798
rect 39849 55795 39915 55798
rect 37273 55722 37339 55725
rect 51625 55722 51691 55725
rect 37273 55720 51691 55722
rect 37273 55664 37278 55720
rect 37334 55664 51630 55720
rect 51686 55664 51691 55720
rect 37273 55662 51691 55664
rect 37273 55659 37339 55662
rect 51625 55659 51691 55662
rect 29269 55586 29335 55589
rect 32857 55586 32923 55589
rect 29269 55584 32923 55586
rect 29269 55528 29274 55584
rect 29330 55528 32862 55584
rect 32918 55528 32923 55584
rect 29269 55526 32923 55528
rect 29269 55523 29335 55526
rect 32857 55523 32923 55526
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 36445 55314 36511 55317
rect 52729 55314 52795 55317
rect 36445 55312 52795 55314
rect 36445 55256 36450 55312
rect 36506 55256 52734 55312
rect 52790 55256 52795 55312
rect 36445 55254 52795 55256
rect 36445 55251 36511 55254
rect 52729 55251 52795 55254
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 24669 2954 24735 2957
rect 31753 2954 31819 2957
rect 24669 2952 31819 2954
rect 24669 2896 24674 2952
rect 24730 2896 31758 2952
rect 31814 2896 31819 2952
rect 24669 2894 31819 2896
rect 24669 2891 24735 2894
rect 31753 2891 31819 2894
rect 35525 2818 35591 2821
rect 38653 2818 38719 2821
rect 35525 2816 38719 2818
rect 35525 2760 35530 2816
rect 35586 2760 38658 2816
rect 38714 2760 38719 2816
rect 35525 2758 38719 2760
rect 35525 2755 35591 2758
rect 38653 2755 38719 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26404 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1666464484
transform 1 0 22080 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1666464484
transform -1 0 31464 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1666464484
transform 1 0 28888 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1666464484
transform 1 0 26312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1666464484
transform 1 0 24012 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A_N
timestamp 1666464484
transform 1 0 36616 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B
timestamp 1666464484
transform 1 0 37076 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__B1
timestamp 1666464484
transform 1 0 29072 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A_N
timestamp 1666464484
transform 1 0 46184 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__B1
timestamp 1666464484
transform 1 0 42228 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B1
timestamp 1666464484
transform -1 0 27416 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1666464484
transform 1 0 34224 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__B2
timestamp 1666464484
transform -1 0 32660 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A2
timestamp 1666464484
transform 1 0 30636 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1666464484
transform 1 0 39560 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A2
timestamp 1666464484
transform -1 0 40848 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1666464484
transform -1 0 23276 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1666464484
transform 1 0 24288 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A2
timestamp 1666464484
transform 1 0 35328 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A2
timestamp 1666464484
transform -1 0 34408 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A1
timestamp 1666464484
transform -1 0 33856 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A1
timestamp 1666464484
transform 1 0 43884 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1666464484
transform 1 0 25116 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1666464484
transform 1 0 24656 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A1
timestamp 1666464484
transform 1 0 33120 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1666464484
transform -1 0 33304 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B1
timestamp 1666464484
transform 1 0 31280 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A1
timestamp 1666464484
transform 1 0 30268 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__B1
timestamp 1666464484
transform 1 0 40756 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A1
timestamp 1666464484
transform 1 0 41308 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A
timestamp 1666464484
transform -1 0 25852 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1666464484
transform 1 0 26496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1666464484
transform 1 0 27416 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A2
timestamp 1666464484
transform 1 0 34776 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A2
timestamp 1666464484
transform -1 0 34960 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A1
timestamp 1666464484
transform -1 0 26772 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__C1
timestamp 1666464484
transform 1 0 28520 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 3864 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 27968 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 24656 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 36248 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 36064 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 35512 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 37444 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 38640 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666464484
transform -1 0 40388 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666464484
transform -1 0 40388 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666464484
transform -1 0 45172 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1666464484
transform -1 0 44620 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1666464484
transform -1 0 46920 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1666464484
transform -1 0 45724 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1666464484
transform -1 0 47472 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1666464484
transform -1 0 48484 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1666464484
transform -1 0 49772 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1666464484
transform -1 0 51428 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1666464484
transform -1 0 52532 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1666464484
transform -1 0 54372 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1666464484
transform -1 0 55844 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output22_A
timestamp 1666464484
transform -1 0 5704 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1666464484
transform 1 0 11040 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33
timestamp 1666464484
transform 1 0 4140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45
timestamp 1666464484
transform 1 0 5244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1666464484
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65
timestamp 1666464484
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1666464484
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1666464484
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87
timestamp 1666464484
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9752 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101
timestamp 1666464484
transform 1 0 10396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_105
timestamp 1666464484
transform 1 0 10764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp 1666464484
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp 1666464484
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129
timestamp 1666464484
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_133
timestamp 1666464484
transform 1 0 13340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144
timestamp 1666464484
transform 1 0 14352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1666464484
transform 1 0 14996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_158
timestamp 1666464484
transform 1 0 15640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_161
timestamp 1666464484
transform 1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_176
timestamp 1666464484
transform 1 0 17296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_183
timestamp 1666464484
transform 1 0 17940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_190
timestamp 1666464484
transform 1 0 18584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_201
timestamp 1666464484
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_208
timestamp 1666464484
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_215
timestamp 1666464484
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1666464484
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_229
timestamp 1666464484
transform 1 0 22172 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1666464484
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1666464484
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1666464484
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_254
timestamp 1666464484
transform 1 0 24472 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_257 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24748 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_286
timestamp 1666464484
transform 1 0 27416 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_289
timestamp 1666464484
transform 1 0 27692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_318
timestamp 1666464484
transform 1 0 30360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp 1666464484
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_344
timestamp 1666464484
transform 1 0 32752 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_353
timestamp 1666464484
transform 1 0 33580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_376
timestamp 1666464484
transform 1 0 35696 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_385
timestamp 1666464484
transform 1 0 36524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_390
timestamp 1666464484
transform 1 0 36984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_397
timestamp 1666464484
transform 1 0 37628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_404
timestamp 1666464484
transform 1 0 38272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_411
timestamp 1666464484
transform 1 0 38916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_415
timestamp 1666464484
transform 1 0 39284 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_417
timestamp 1666464484
transform 1 0 39468 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_422
timestamp 1666464484
transform 1 0 39928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1666464484
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_436
timestamp 1666464484
transform 1 0 41216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_443
timestamp 1666464484
transform 1 0 41860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1666464484
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1666464484
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_454
timestamp 1666464484
transform 1 0 42872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1666464484
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_468
timestamp 1666464484
transform 1 0 44160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_475
timestamp 1666464484
transform 1 0 44804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_479
timestamp 1666464484
transform 1 0 45172 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_481
timestamp 1666464484
transform 1 0 45356 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_486
timestamp 1666464484
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_493
timestamp 1666464484
transform 1 0 46460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1666464484
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_507
timestamp 1666464484
transform 1 0 47748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_511
timestamp 1666464484
transform 1 0 48116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_513
timestamp 1666464484
transform 1 0 48300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_518
timestamp 1666464484
transform 1 0 48760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_525
timestamp 1666464484
transform 1 0 49404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_532
timestamp 1666464484
transform 1 0 50048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_539
timestamp 1666464484
transform 1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_543
timestamp 1666464484
transform 1 0 51060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_545
timestamp 1666464484
transform 1 0 51244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_550
timestamp 1666464484
transform 1 0 51704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_557
timestamp 1666464484
transform 1 0 52348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_564
timestamp 1666464484
transform 1 0 52992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_571
timestamp 1666464484
transform 1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_575
timestamp 1666464484
transform 1 0 54004 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_577
timestamp 1666464484
transform 1 0 54188 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1666464484
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_601
timestamp 1666464484
transform 1 0 56396 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_607
timestamp 1666464484
transform 1 0 56948 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_609
timestamp 1666464484
transform 1 0 57132 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_621
timestamp 1666464484
transform 1 0 58236 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_51
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_63
timestamp 1666464484
transform 1 0 6900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_66
timestamp 1666464484
transform 1 0 7176 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_75
timestamp 1666464484
transform 1 0 8004 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85
timestamp 1666464484
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_89
timestamp 1666464484
transform 1 0 9292 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_100
timestamp 1666464484
transform 1 0 10304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1666464484
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_114
timestamp 1666464484
transform 1 0 11592 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_121
timestamp 1666464484
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_128
timestamp 1666464484
transform 1 0 12880 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_131 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_144
timestamp 1666464484
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_151
timestamp 1666464484
transform 1 0 14996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp 1666464484
transform 1 0 15640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_165
timestamp 1666464484
transform 1 0 16284 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1666464484
transform 1 0 16928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1666464484
transform 1 0 17572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_186
timestamp 1666464484
transform 1 0 18216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_196
timestamp 1666464484
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1666464484
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp 1666464484
transform 1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_216
timestamp 1666464484
transform 1 0 20976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_230
timestamp 1666464484
transform 1 0 22264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1666464484
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1666464484
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_251
timestamp 1666464484
transform 1 0 24196 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_258
timestamp 1666464484
transform 1 0 24840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_261
timestamp 1666464484
transform 1 0 25116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_265
timestamp 1666464484
transform 1 0 25484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_287
timestamp 1666464484
transform 1 0 27508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_312
timestamp 1666464484
transform 1 0 29808 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_323
timestamp 1666464484
transform 1 0 30820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_326
timestamp 1666464484
transform 1 0 31096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_330
timestamp 1666464484
transform 1 0 31464 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_352
timestamp 1666464484
transform 1 0 33488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_377
timestamp 1666464484
transform 1 0 35788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_384
timestamp 1666464484
transform 1 0 36432 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_391
timestamp 1666464484
transform 1 0 37076 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_396
timestamp 1666464484
transform 1 0 37536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1666464484
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_410
timestamp 1666464484
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1666464484
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1666464484
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1666464484
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_438
timestamp 1666464484
transform 1 0 41400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_445
timestamp 1666464484
transform 1 0 42044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_452
timestamp 1666464484
transform 1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_456
timestamp 1666464484
transform 1 0 43056 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1666464484
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_468
timestamp 1666464484
transform 1 0 44160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_475
timestamp 1666464484
transform 1 0 44804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1666464484
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_489
timestamp 1666464484
transform 1 0 46092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_496
timestamp 1666464484
transform 1 0 46736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_503
timestamp 1666464484
transform 1 0 47380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_510
timestamp 1666464484
transform 1 0 48024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_517
timestamp 1666464484
transform 1 0 48668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_521
timestamp 1666464484
transform 1 0 49036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_526
timestamp 1666464484
transform 1 0 49496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_533
timestamp 1666464484
transform 1 0 50140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_540
timestamp 1666464484
transform 1 0 50784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_547
timestamp 1666464484
transform 1 0 51428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_554
timestamp 1666464484
transform 1 0 52072 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_561
timestamp 1666464484
transform 1 0 52716 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_568
timestamp 1666464484
transform 1 0 53360 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_580
timestamp 1666464484
transform 1 0 54464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_584
timestamp 1666464484
transform 1 0 54832 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_586
timestamp 1666464484
transform 1 0 55016 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_598
timestamp 1666464484
transform 1 0 56120 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_610
timestamp 1666464484
transform 1 0 57224 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_622
timestamp 1666464484
transform 1 0 58328 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_31
timestamp 1666464484
transform 1 0 3956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_33
timestamp 1666464484
transform 1 0 4140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_45
timestamp 1666464484
transform 1 0 5244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_57
timestamp 1666464484
transform 1 0 6348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_69
timestamp 1666464484
transform 1 0 7452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_81
timestamp 1666464484
transform 1 0 8556 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1666464484
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1666464484
transform 1 0 9660 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_98
timestamp 1666464484
transform 1 0 10120 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_127
timestamp 1666464484
transform 1 0 12788 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_135
timestamp 1666464484
transform 1 0 13524 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_147
timestamp 1666464484
transform 1 0 14628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_151
timestamp 1666464484
transform 1 0 14996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_160
timestamp 1666464484
transform 1 0 15824 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_163
timestamp 1666464484
transform 1 0 16100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1666464484
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_176
timestamp 1666464484
transform 1 0 17296 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_180
timestamp 1666464484
transform 1 0 17664 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_193
timestamp 1666464484
transform 1 0 18860 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_204
timestamp 1666464484
transform 1 0 19872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_211
timestamp 1666464484
transform 1 0 20516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_218
timestamp 1666464484
transform 1 0 21160 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_225
timestamp 1666464484
transform 1 0 21804 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_228
timestamp 1666464484
transform 1 0 22080 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_233
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1666464484
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_265
timestamp 1666464484
transform 1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_290
timestamp 1666464484
transform 1 0 27784 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_293
timestamp 1666464484
transform 1 0 28060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_316
timestamp 1666464484
transform 1 0 30176 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_325
timestamp 1666464484
transform 1 0 31004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_329
timestamp 1666464484
transform 1 0 31372 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_351
timestamp 1666464484
transform 1 0 33396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_358
timestamp 1666464484
transform 1 0 34040 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_381
timestamp 1666464484
transform 1 0 36156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_388
timestamp 1666464484
transform 1 0 36800 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_395
timestamp 1666464484
transform 1 0 37444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_402
timestamp 1666464484
transform 1 0 38088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_409
timestamp 1666464484
transform 1 0 38732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_416
timestamp 1666464484
transform 1 0 39376 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_423
timestamp 1666464484
transform 1 0 40020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_428
timestamp 1666464484
transform 1 0 40480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_435
timestamp 1666464484
transform 1 0 41124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_442
timestamp 1666464484
transform 1 0 41768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_449
timestamp 1666464484
transform 1 0 42412 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_456
timestamp 1666464484
transform 1 0 43056 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_463
timestamp 1666464484
transform 1 0 43700 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_467
timestamp 1666464484
transform 1 0 44068 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_471
timestamp 1666464484
transform 1 0 44436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_483
timestamp 1666464484
transform 1 0 45540 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_488
timestamp 1666464484
transform 1 0 46000 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_493
timestamp 1666464484
transform 1 0 46460 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_500
timestamp 1666464484
transform 1 0 47104 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_512
timestamp 1666464484
transform 1 0 48208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_516
timestamp 1666464484
transform 1 0 48576 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_524
timestamp 1666464484
transform 1 0 49312 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_528
timestamp 1666464484
transform 1 0 49680 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_537
timestamp 1666464484
transform 1 0 50508 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_549
timestamp 1666464484
transform 1 0 51612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_553
timestamp 1666464484
transform 1 0 51980 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_558
timestamp 1666464484
transform 1 0 52440 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_570
timestamp 1666464484
transform 1 0 53544 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_582
timestamp 1666464484
transform 1 0 54648 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_594
timestamp 1666464484
transform 1 0 55752 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_606
timestamp 1666464484
transform 1 0 56856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_614
timestamp 1666464484
transform 1 0 57592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_618
timestamp 1666464484
transform 1 0 57960 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_624
timestamp 1666464484
transform 1 0 58512 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666464484
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_51
timestamp 1666464484
transform 1 0 5796 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_63
timestamp 1666464484
transform 1 0 6900 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_66
timestamp 1666464484
transform 1 0 7176 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_78
timestamp 1666464484
transform 1 0 8280 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_90
timestamp 1666464484
transform 1 0 9384 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_102
timestamp 1666464484
transform 1 0 10488 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_114
timestamp 1666464484
transform 1 0 11592 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_126
timestamp 1666464484
transform 1 0 12696 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_131
timestamp 1666464484
transform 1 0 13156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_143
timestamp 1666464484
transform 1 0 14260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_155
timestamp 1666464484
transform 1 0 15364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_179
timestamp 1666464484
transform 1 0 17572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_191
timestamp 1666464484
transform 1 0 18676 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_196
timestamp 1666464484
transform 1 0 19136 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_207
timestamp 1666464484
transform 1 0 20148 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_216
timestamp 1666464484
transform 1 0 20976 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_223
timestamp 1666464484
transform 1 0 21620 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_230
timestamp 1666464484
transform 1 0 22264 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_237
timestamp 1666464484
transform 1 0 22908 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1666464484
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_251
timestamp 1666464484
transform 1 0 24196 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_258
timestamp 1666464484
transform 1 0 24840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_261
timestamp 1666464484
transform 1 0 25116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_266
timestamp 1666464484
transform 1 0 25576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_273
timestamp 1666464484
transform 1 0 26220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_298
timestamp 1666464484
transform 1 0 28520 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_323
timestamp 1666464484
transform 1 0 30820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_326
timestamp 1666464484
transform 1 0 31096 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_331
timestamp 1666464484
transform 1 0 31556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_338
timestamp 1666464484
transform 1 0 32200 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_342
timestamp 1666464484
transform 1 0 32568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_364
timestamp 1666464484
transform 1 0 34592 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_371
timestamp 1666464484
transform 1 0 35236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_378
timestamp 1666464484
transform 1 0 35880 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_385
timestamp 1666464484
transform 1 0 36524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_389
timestamp 1666464484
transform 1 0 36892 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_391
timestamp 1666464484
transform 1 0 37076 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_396
timestamp 1666464484
transform 1 0 37536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1666464484
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_407
timestamp 1666464484
transform 1 0 38548 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_411
timestamp 1666464484
transform 1 0 38916 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_423
timestamp 1666464484
transform 1 0 40020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_435
timestamp 1666464484
transform 1 0 41124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_447
timestamp 1666464484
transform 1 0 42228 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_456
timestamp 1666464484
transform 1 0 43056 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_468
timestamp 1666464484
transform 1 0 44160 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_480
timestamp 1666464484
transform 1 0 45264 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_492
timestamp 1666464484
transform 1 0 46368 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_504
timestamp 1666464484
transform 1 0 47472 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_516
timestamp 1666464484
transform 1 0 48576 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_521
timestamp 1666464484
transform 1 0 49036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_533
timestamp 1666464484
transform 1 0 50140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_545
timestamp 1666464484
transform 1 0 51244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_557
timestamp 1666464484
transform 1 0 52348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_569
timestamp 1666464484
transform 1 0 53452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_581
timestamp 1666464484
transform 1 0 54556 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_586
timestamp 1666464484
transform 1 0 55016 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_598
timestamp 1666464484
transform 1 0 56120 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_610
timestamp 1666464484
transform 1 0 57224 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_622
timestamp 1666464484
transform 1 0 58328 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_31
timestamp 1666464484
transform 1 0 3956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_33
timestamp 1666464484
transform 1 0 4140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_45
timestamp 1666464484
transform 1 0 5244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_57
timestamp 1666464484
transform 1 0 6348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_69
timestamp 1666464484
transform 1 0 7452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_81
timestamp 1666464484
transform 1 0 8556 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1666464484
transform 1 0 9660 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_98
timestamp 1666464484
transform 1 0 10120 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_110
timestamp 1666464484
transform 1 0 11224 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_122
timestamp 1666464484
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_134
timestamp 1666464484
transform 1 0 13432 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_146
timestamp 1666464484
transform 1 0 14536 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_158
timestamp 1666464484
transform 1 0 15640 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_163
timestamp 1666464484
transform 1 0 16100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_175
timestamp 1666464484
transform 1 0 17204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_187
timestamp 1666464484
transform 1 0 18308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_199
timestamp 1666464484
transform 1 0 19412 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_211
timestamp 1666464484
transform 1 0 20516 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_219
timestamp 1666464484
transform 1 0 21252 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_225
timestamp 1666464484
transform 1 0 21804 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_228
timestamp 1666464484
transform 1 0 22080 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_237
timestamp 1666464484
transform 1 0 22908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_244
timestamp 1666464484
transform 1 0 23552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_251
timestamp 1666464484
transform 1 0 24196 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_258
timestamp 1666464484
transform 1 0 24840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_290
timestamp 1666464484
transform 1 0 27784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_293
timestamp 1666464484
transform 1 0 28060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_299
timestamp 1666464484
transform 1 0 28612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_306
timestamp 1666464484
transform 1 0 29256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_313
timestamp 1666464484
transform 1 0 29900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_338
timestamp 1666464484
transform 1 0 32200 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_345
timestamp 1666464484
transform 1 0 32844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_352
timestamp 1666464484
transform 1 0 33488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_356
timestamp 1666464484
transform 1 0 33856 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_358
timestamp 1666464484
transform 1 0 34040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_381
timestamp 1666464484
transform 1 0 36156 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_388
timestamp 1666464484
transform 1 0 36800 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_400
timestamp 1666464484
transform 1 0 37904 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_412
timestamp 1666464484
transform 1 0 39008 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_420
timestamp 1666464484
transform 1 0 39744 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_423
timestamp 1666464484
transform 1 0 40020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_435
timestamp 1666464484
transform 1 0 41124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_447
timestamp 1666464484
transform 1 0 42228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_459
timestamp 1666464484
transform 1 0 43332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_471
timestamp 1666464484
transform 1 0 44436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_483
timestamp 1666464484
transform 1 0 45540 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_488
timestamp 1666464484
transform 1 0 46000 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_500
timestamp 1666464484
transform 1 0 47104 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_512
timestamp 1666464484
transform 1 0 48208 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_524
timestamp 1666464484
transform 1 0 49312 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_536
timestamp 1666464484
transform 1 0 50416 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_548
timestamp 1666464484
transform 1 0 51520 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_553
timestamp 1666464484
transform 1 0 51980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_565
timestamp 1666464484
transform 1 0 53084 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_577
timestamp 1666464484
transform 1 0 54188 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1666464484
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1666464484
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_613
timestamp 1666464484
transform 1 0 57500 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_618
timestamp 1666464484
transform 1 0 57960 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_624
timestamp 1666464484
transform 1 0 58512 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1666464484
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_51
timestamp 1666464484
transform 1 0 5796 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_63
timestamp 1666464484
transform 1 0 6900 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_66
timestamp 1666464484
transform 1 0 7176 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_78
timestamp 1666464484
transform 1 0 8280 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_90
timestamp 1666464484
transform 1 0 9384 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_102
timestamp 1666464484
transform 1 0 10488 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_114
timestamp 1666464484
transform 1 0 11592 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_126
timestamp 1666464484
transform 1 0 12696 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_131
timestamp 1666464484
transform 1 0 13156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_143
timestamp 1666464484
transform 1 0 14260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_155
timestamp 1666464484
transform 1 0 15364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_179
timestamp 1666464484
transform 1 0 17572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1666464484
transform 1 0 18676 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_196
timestamp 1666464484
transform 1 0 19136 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_208
timestamp 1666464484
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_220
timestamp 1666464484
transform 1 0 21344 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_232
timestamp 1666464484
transform 1 0 22448 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1666464484
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1666464484
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_251
timestamp 1666464484
transform 1 0 24196 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_258
timestamp 1666464484
transform 1 0 24840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_284
timestamp 1666464484
transform 1 0 27232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_291
timestamp 1666464484
transform 1 0 27876 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_298
timestamp 1666464484
transform 1 0 28520 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_323
timestamp 1666464484
transform 1 0 30820 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_326
timestamp 1666464484
transform 1 0 31096 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_349
timestamp 1666464484
transform 1 0 33212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_374
timestamp 1666464484
transform 1 0 35512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_381
timestamp 1666464484
transform 1 0 36156 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_389
timestamp 1666464484
transform 1 0 36892 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_391
timestamp 1666464484
transform 1 0 37076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_403
timestamp 1666464484
transform 1 0 38180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_415
timestamp 1666464484
transform 1 0 39284 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_427
timestamp 1666464484
transform 1 0 40388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_439
timestamp 1666464484
transform 1 0 41492 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_451
timestamp 1666464484
transform 1 0 42596 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_456
timestamp 1666464484
transform 1 0 43056 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_468
timestamp 1666464484
transform 1 0 44160 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_480
timestamp 1666464484
transform 1 0 45264 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_492
timestamp 1666464484
transform 1 0 46368 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_504
timestamp 1666464484
transform 1 0 47472 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_516
timestamp 1666464484
transform 1 0 48576 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_521
timestamp 1666464484
transform 1 0 49036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_533
timestamp 1666464484
transform 1 0 50140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_545
timestamp 1666464484
transform 1 0 51244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_557
timestamp 1666464484
transform 1 0 52348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_569
timestamp 1666464484
transform 1 0 53452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_581
timestamp 1666464484
transform 1 0 54556 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_586
timestamp 1666464484
transform 1 0 55016 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_598
timestamp 1666464484
transform 1 0 56120 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_610
timestamp 1666464484
transform 1 0 57224 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_622
timestamp 1666464484
transform 1 0 58328 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_31
timestamp 1666464484
transform 1 0 3956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_33
timestamp 1666464484
transform 1 0 4140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_45
timestamp 1666464484
transform 1 0 5244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_57
timestamp 1666464484
transform 1 0 6348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_69
timestamp 1666464484
transform 1 0 7452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_81
timestamp 1666464484
transform 1 0 8556 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1666464484
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_98
timestamp 1666464484
transform 1 0 10120 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_110
timestamp 1666464484
transform 1 0 11224 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_122
timestamp 1666464484
transform 1 0 12328 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_134
timestamp 1666464484
transform 1 0 13432 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_146
timestamp 1666464484
transform 1 0 14536 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_158
timestamp 1666464484
transform 1 0 15640 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_163
timestamp 1666464484
transform 1 0 16100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_175
timestamp 1666464484
transform 1 0 17204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_187
timestamp 1666464484
transform 1 0 18308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_199
timestamp 1666464484
transform 1 0 19412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_211
timestamp 1666464484
transform 1 0 20516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1666464484
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_228
timestamp 1666464484
transform 1 0 22080 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_240
timestamp 1666464484
transform 1 0 23184 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_248
timestamp 1666464484
transform 1 0 23920 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_258
timestamp 1666464484
transform 1 0 24840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_290
timestamp 1666464484
transform 1 0 27784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_293
timestamp 1666464484
transform 1 0 28060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_299
timestamp 1666464484
transform 1 0 28612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1666464484
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_310
timestamp 1666464484
transform 1 0 29624 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_335
timestamp 1666464484
transform 1 0 31924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_342
timestamp 1666464484
transform 1 0 32568 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_349
timestamp 1666464484
transform 1 0 33212 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_358
timestamp 1666464484
transform 1 0 34040 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_381
timestamp 1666464484
transform 1 0 36156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_393
timestamp 1666464484
transform 1 0 37260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_405
timestamp 1666464484
transform 1 0 38364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_417
timestamp 1666464484
transform 1 0 39468 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_421
timestamp 1666464484
transform 1 0 39836 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_423
timestamp 1666464484
transform 1 0 40020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_435
timestamp 1666464484
transform 1 0 41124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_447
timestamp 1666464484
transform 1 0 42228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_459
timestamp 1666464484
transform 1 0 43332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_471
timestamp 1666464484
transform 1 0 44436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_483
timestamp 1666464484
transform 1 0 45540 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_488
timestamp 1666464484
transform 1 0 46000 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_500
timestamp 1666464484
transform 1 0 47104 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_512
timestamp 1666464484
transform 1 0 48208 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_524
timestamp 1666464484
transform 1 0 49312 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_536
timestamp 1666464484
transform 1 0 50416 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_548
timestamp 1666464484
transform 1 0 51520 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_553
timestamp 1666464484
transform 1 0 51980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_565
timestamp 1666464484
transform 1 0 53084 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_577
timestamp 1666464484
transform 1 0 54188 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1666464484
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1666464484
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_613
timestamp 1666464484
transform 1 0 57500 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_618
timestamp 1666464484
transform 1 0 57960 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_624
timestamp 1666464484
transform 1 0 58512 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_51
timestamp 1666464484
transform 1 0 5796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_63
timestamp 1666464484
transform 1 0 6900 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_66
timestamp 1666464484
transform 1 0 7176 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_78
timestamp 1666464484
transform 1 0 8280 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_90
timestamp 1666464484
transform 1 0 9384 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_102
timestamp 1666464484
transform 1 0 10488 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_114
timestamp 1666464484
transform 1 0 11592 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_126
timestamp 1666464484
transform 1 0 12696 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_131
timestamp 1666464484
transform 1 0 13156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_143
timestamp 1666464484
transform 1 0 14260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_155
timestamp 1666464484
transform 1 0 15364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_179
timestamp 1666464484
transform 1 0 17572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp 1666464484
transform 1 0 18676 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_196
timestamp 1666464484
transform 1 0 19136 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_208
timestamp 1666464484
transform 1 0 20240 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_220
timestamp 1666464484
transform 1 0 21344 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_232
timestamp 1666464484
transform 1 0 22448 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_244
timestamp 1666464484
transform 1 0 23552 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_256
timestamp 1666464484
transform 1 0 24656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_266
timestamp 1666464484
transform 1 0 25576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_270
timestamp 1666464484
transform 1 0 25944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_274
timestamp 1666464484
transform 1 0 26312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_284
timestamp 1666464484
transform 1 0 27232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_309
timestamp 1666464484
transform 1 0 29532 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_323
timestamp 1666464484
transform 1 0 30820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_326
timestamp 1666464484
transform 1 0 31096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_330
timestamp 1666464484
transform 1 0 31464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_355
timestamp 1666464484
transform 1 0 33764 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_362
timestamp 1666464484
transform 1 0 34408 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_374
timestamp 1666464484
transform 1 0 35512 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_386
timestamp 1666464484
transform 1 0 36616 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_391
timestamp 1666464484
transform 1 0 37076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_403
timestamp 1666464484
transform 1 0 38180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_415
timestamp 1666464484
transform 1 0 39284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_427
timestamp 1666464484
transform 1 0 40388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_439
timestamp 1666464484
transform 1 0 41492 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_451
timestamp 1666464484
transform 1 0 42596 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_456
timestamp 1666464484
transform 1 0 43056 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_468
timestamp 1666464484
transform 1 0 44160 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_480
timestamp 1666464484
transform 1 0 45264 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_492
timestamp 1666464484
transform 1 0 46368 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_504
timestamp 1666464484
transform 1 0 47472 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_516
timestamp 1666464484
transform 1 0 48576 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_521
timestamp 1666464484
transform 1 0 49036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_533
timestamp 1666464484
transform 1 0 50140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_545
timestamp 1666464484
transform 1 0 51244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_557
timestamp 1666464484
transform 1 0 52348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_569
timestamp 1666464484
transform 1 0 53452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_581
timestamp 1666464484
transform 1 0 54556 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_586
timestamp 1666464484
transform 1 0 55016 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_598
timestamp 1666464484
transform 1 0 56120 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_610
timestamp 1666464484
transform 1 0 57224 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_622
timestamp 1666464484
transform 1 0 58328 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_31
timestamp 1666464484
transform 1 0 3956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_33
timestamp 1666464484
transform 1 0 4140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_45
timestamp 1666464484
transform 1 0 5244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_57
timestamp 1666464484
transform 1 0 6348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_69
timestamp 1666464484
transform 1 0 7452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_81
timestamp 1666464484
transform 1 0 8556 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1666464484
transform 1 0 9660 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_98
timestamp 1666464484
transform 1 0 10120 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_110
timestamp 1666464484
transform 1 0 11224 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_122
timestamp 1666464484
transform 1 0 12328 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_134
timestamp 1666464484
transform 1 0 13432 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_146
timestamp 1666464484
transform 1 0 14536 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_158
timestamp 1666464484
transform 1 0 15640 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_163
timestamp 1666464484
transform 1 0 16100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_175
timestamp 1666464484
transform 1 0 17204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_187
timestamp 1666464484
transform 1 0 18308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_199
timestamp 1666464484
transform 1 0 19412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_211
timestamp 1666464484
transform 1 0 20516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_223
timestamp 1666464484
transform 1 0 21620 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_228
timestamp 1666464484
transform 1 0 22080 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_240
timestamp 1666464484
transform 1 0 23184 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_252
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_264
timestamp 1666464484
transform 1 0 25392 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_272
timestamp 1666464484
transform 1 0 26128 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_276
timestamp 1666464484
transform 1 0 26496 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_283
timestamp 1666464484
transform 1 0 27140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_290
timestamp 1666464484
transform 1 0 27784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_293
timestamp 1666464484
transform 1 0 28060 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_299
timestamp 1666464484
transform 1 0 28612 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_321
timestamp 1666464484
transform 1 0 30636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_346
timestamp 1666464484
transform 1 0 32936 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_354
timestamp 1666464484
transform 1 0 33672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_358
timestamp 1666464484
transform 1 0 34040 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_363
timestamp 1666464484
transform 1 0 34500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_375
timestamp 1666464484
transform 1 0 35604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_387
timestamp 1666464484
transform 1 0 36708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_399
timestamp 1666464484
transform 1 0 37812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_411
timestamp 1666464484
transform 1 0 38916 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_419
timestamp 1666464484
transform 1 0 39652 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_423
timestamp 1666464484
transform 1 0 40020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_435
timestamp 1666464484
transform 1 0 41124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_447
timestamp 1666464484
transform 1 0 42228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_459
timestamp 1666464484
transform 1 0 43332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_471
timestamp 1666464484
transform 1 0 44436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_483
timestamp 1666464484
transform 1 0 45540 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_488
timestamp 1666464484
transform 1 0 46000 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_500
timestamp 1666464484
transform 1 0 47104 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_512
timestamp 1666464484
transform 1 0 48208 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_524
timestamp 1666464484
transform 1 0 49312 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_536
timestamp 1666464484
transform 1 0 50416 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_548
timestamp 1666464484
transform 1 0 51520 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_553
timestamp 1666464484
transform 1 0 51980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_565
timestamp 1666464484
transform 1 0 53084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_577
timestamp 1666464484
transform 1 0 54188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1666464484
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1666464484
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_613
timestamp 1666464484
transform 1 0 57500 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_618
timestamp 1666464484
transform 1 0 57960 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_624
timestamp 1666464484
transform 1 0 58512 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666464484
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_51
timestamp 1666464484
transform 1 0 5796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_63
timestamp 1666464484
transform 1 0 6900 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_66
timestamp 1666464484
transform 1 0 7176 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_78
timestamp 1666464484
transform 1 0 8280 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_90
timestamp 1666464484
transform 1 0 9384 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_102
timestamp 1666464484
transform 1 0 10488 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_114
timestamp 1666464484
transform 1 0 11592 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_126
timestamp 1666464484
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_131
timestamp 1666464484
transform 1 0 13156 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_143
timestamp 1666464484
transform 1 0 14260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_155
timestamp 1666464484
transform 1 0 15364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_179
timestamp 1666464484
transform 1 0 17572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_191
timestamp 1666464484
transform 1 0 18676 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_196
timestamp 1666464484
transform 1 0 19136 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_208
timestamp 1666464484
transform 1 0 20240 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_220
timestamp 1666464484
transform 1 0 21344 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_232
timestamp 1666464484
transform 1 0 22448 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_244
timestamp 1666464484
transform 1 0 23552 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_256
timestamp 1666464484
transform 1 0 24656 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1666464484
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1666464484
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_282
timestamp 1666464484
transform 1 0 27048 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_288
timestamp 1666464484
transform 1 0 27600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_310
timestamp 1666464484
transform 1 0 29624 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_320
timestamp 1666464484
transform 1 0 30544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_324
timestamp 1666464484
transform 1 0 30912 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_326
timestamp 1666464484
transform 1 0 31096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_331
timestamp 1666464484
transform 1 0 31556 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_340
timestamp 1666464484
transform 1 0 32384 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_352
timestamp 1666464484
transform 1 0 33488 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_364
timestamp 1666464484
transform 1 0 34592 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_376
timestamp 1666464484
transform 1 0 35696 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_388
timestamp 1666464484
transform 1 0 36800 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_391
timestamp 1666464484
transform 1 0 37076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_403
timestamp 1666464484
transform 1 0 38180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_415
timestamp 1666464484
transform 1 0 39284 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_427
timestamp 1666464484
transform 1 0 40388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_439
timestamp 1666464484
transform 1 0 41492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_451
timestamp 1666464484
transform 1 0 42596 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_456
timestamp 1666464484
transform 1 0 43056 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_468
timestamp 1666464484
transform 1 0 44160 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_480
timestamp 1666464484
transform 1 0 45264 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_492
timestamp 1666464484
transform 1 0 46368 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_504
timestamp 1666464484
transform 1 0 47472 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_516
timestamp 1666464484
transform 1 0 48576 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_521
timestamp 1666464484
transform 1 0 49036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_533
timestamp 1666464484
transform 1 0 50140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_545
timestamp 1666464484
transform 1 0 51244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_557
timestamp 1666464484
transform 1 0 52348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_569
timestamp 1666464484
transform 1 0 53452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_581
timestamp 1666464484
transform 1 0 54556 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_586
timestamp 1666464484
transform 1 0 55016 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_598
timestamp 1666464484
transform 1 0 56120 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_610
timestamp 1666464484
transform 1 0 57224 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_622
timestamp 1666464484
transform 1 0 58328 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_31
timestamp 1666464484
transform 1 0 3956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_33
timestamp 1666464484
transform 1 0 4140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_45
timestamp 1666464484
transform 1 0 5244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_57
timestamp 1666464484
transform 1 0 6348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_69
timestamp 1666464484
transform 1 0 7452 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_81
timestamp 1666464484
transform 1 0 8556 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1666464484
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_98
timestamp 1666464484
transform 1 0 10120 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_110
timestamp 1666464484
transform 1 0 11224 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_122
timestamp 1666464484
transform 1 0 12328 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_134
timestamp 1666464484
transform 1 0 13432 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_146
timestamp 1666464484
transform 1 0 14536 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_158
timestamp 1666464484
transform 1 0 15640 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_163
timestamp 1666464484
transform 1 0 16100 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_175
timestamp 1666464484
transform 1 0 17204 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_187
timestamp 1666464484
transform 1 0 18308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_199
timestamp 1666464484
transform 1 0 19412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_211
timestamp 1666464484
transform 1 0 20516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1666464484
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_228
timestamp 1666464484
transform 1 0 22080 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_240
timestamp 1666464484
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_252
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_264
timestamp 1666464484
transform 1 0 25392 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_276
timestamp 1666464484
transform 1 0 26496 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_288
timestamp 1666464484
transform 1 0 27600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_293
timestamp 1666464484
transform 1 0 28060 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_301
timestamp 1666464484
transform 1 0 28796 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1666464484
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_311
timestamp 1666464484
transform 1 0 29716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_318
timestamp 1666464484
transform 1 0 30360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_322
timestamp 1666464484
transform 1 0 30728 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_326
timestamp 1666464484
transform 1 0 31096 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_338
timestamp 1666464484
transform 1 0 32200 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_350
timestamp 1666464484
transform 1 0 33304 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_356
timestamp 1666464484
transform 1 0 33856 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_358
timestamp 1666464484
transform 1 0 34040 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_370
timestamp 1666464484
transform 1 0 35144 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_382
timestamp 1666464484
transform 1 0 36248 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_394
timestamp 1666464484
transform 1 0 37352 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_406
timestamp 1666464484
transform 1 0 38456 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_418
timestamp 1666464484
transform 1 0 39560 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_423
timestamp 1666464484
transform 1 0 40020 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_435
timestamp 1666464484
transform 1 0 41124 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_447
timestamp 1666464484
transform 1 0 42228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_459
timestamp 1666464484
transform 1 0 43332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_471
timestamp 1666464484
transform 1 0 44436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_483
timestamp 1666464484
transform 1 0 45540 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_488
timestamp 1666464484
transform 1 0 46000 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_500
timestamp 1666464484
transform 1 0 47104 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_512
timestamp 1666464484
transform 1 0 48208 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_524
timestamp 1666464484
transform 1 0 49312 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_536
timestamp 1666464484
transform 1 0 50416 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_548
timestamp 1666464484
transform 1 0 51520 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_553
timestamp 1666464484
transform 1 0 51980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_565
timestamp 1666464484
transform 1 0 53084 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_577
timestamp 1666464484
transform 1 0 54188 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1666464484
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1666464484
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_613
timestamp 1666464484
transform 1 0 57500 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_618
timestamp 1666464484
transform 1 0 57960 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_624
timestamp 1666464484
transform 1 0 58512 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_63
timestamp 1666464484
transform 1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_66
timestamp 1666464484
transform 1 0 7176 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_78
timestamp 1666464484
transform 1 0 8280 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_90
timestamp 1666464484
transform 1 0 9384 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_102
timestamp 1666464484
transform 1 0 10488 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_114
timestamp 1666464484
transform 1 0 11592 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_126
timestamp 1666464484
transform 1 0 12696 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_131
timestamp 1666464484
transform 1 0 13156 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_143
timestamp 1666464484
transform 1 0 14260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_155
timestamp 1666464484
transform 1 0 15364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_179
timestamp 1666464484
transform 1 0 17572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1666464484
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_196
timestamp 1666464484
transform 1 0 19136 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_208
timestamp 1666464484
transform 1 0 20240 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_220
timestamp 1666464484
transform 1 0 21344 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_232
timestamp 1666464484
transform 1 0 22448 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_244
timestamp 1666464484
transform 1 0 23552 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_256
timestamp 1666464484
transform 1 0 24656 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1666464484
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_273
timestamp 1666464484
transform 1 0 26220 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_285
timestamp 1666464484
transform 1 0 27324 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_297
timestamp 1666464484
transform 1 0 28428 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_309
timestamp 1666464484
transform 1 0 29532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_313
timestamp 1666464484
transform 1 0 29900 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_317
timestamp 1666464484
transform 1 0 30268 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_326
timestamp 1666464484
transform 1 0 31096 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_338
timestamp 1666464484
transform 1 0 32200 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_350
timestamp 1666464484
transform 1 0 33304 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_362
timestamp 1666464484
transform 1 0 34408 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_374
timestamp 1666464484
transform 1 0 35512 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_386
timestamp 1666464484
transform 1 0 36616 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_391
timestamp 1666464484
transform 1 0 37076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_403
timestamp 1666464484
transform 1 0 38180 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_415
timestamp 1666464484
transform 1 0 39284 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_427
timestamp 1666464484
transform 1 0 40388 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_439
timestamp 1666464484
transform 1 0 41492 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_451
timestamp 1666464484
transform 1 0 42596 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_456
timestamp 1666464484
transform 1 0 43056 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_468
timestamp 1666464484
transform 1 0 44160 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_480
timestamp 1666464484
transform 1 0 45264 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_492
timestamp 1666464484
transform 1 0 46368 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_504
timestamp 1666464484
transform 1 0 47472 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_516
timestamp 1666464484
transform 1 0 48576 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_521
timestamp 1666464484
transform 1 0 49036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_533
timestamp 1666464484
transform 1 0 50140 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_545
timestamp 1666464484
transform 1 0 51244 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_557
timestamp 1666464484
transform 1 0 52348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_569
timestamp 1666464484
transform 1 0 53452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_581
timestamp 1666464484
transform 1 0 54556 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_586
timestamp 1666464484
transform 1 0 55016 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_598
timestamp 1666464484
transform 1 0 56120 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_610
timestamp 1666464484
transform 1 0 57224 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_622
timestamp 1666464484
transform 1 0 58328 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_31
timestamp 1666464484
transform 1 0 3956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_33
timestamp 1666464484
transform 1 0 4140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_45
timestamp 1666464484
transform 1 0 5244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_57
timestamp 1666464484
transform 1 0 6348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_69
timestamp 1666464484
transform 1 0 7452 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_81
timestamp 1666464484
transform 1 0 8556 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1666464484
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_98
timestamp 1666464484
transform 1 0 10120 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_110
timestamp 1666464484
transform 1 0 11224 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_122
timestamp 1666464484
transform 1 0 12328 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_134
timestamp 1666464484
transform 1 0 13432 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_146
timestamp 1666464484
transform 1 0 14536 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_158
timestamp 1666464484
transform 1 0 15640 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_163
timestamp 1666464484
transform 1 0 16100 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_175
timestamp 1666464484
transform 1 0 17204 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_187
timestamp 1666464484
transform 1 0 18308 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_199
timestamp 1666464484
transform 1 0 19412 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_211
timestamp 1666464484
transform 1 0 20516 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_223
timestamp 1666464484
transform 1 0 21620 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_228
timestamp 1666464484
transform 1 0 22080 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_240
timestamp 1666464484
transform 1 0 23184 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_252
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_264
timestamp 1666464484
transform 1 0 25392 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_276
timestamp 1666464484
transform 1 0 26496 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_288
timestamp 1666464484
transform 1 0 27600 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_293
timestamp 1666464484
transform 1 0 28060 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_305
timestamp 1666464484
transform 1 0 29164 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_317
timestamp 1666464484
transform 1 0 30268 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_329
timestamp 1666464484
transform 1 0 31372 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_341
timestamp 1666464484
transform 1 0 32476 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_353
timestamp 1666464484
transform 1 0 33580 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_358
timestamp 1666464484
transform 1 0 34040 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_370
timestamp 1666464484
transform 1 0 35144 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_382
timestamp 1666464484
transform 1 0 36248 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_394
timestamp 1666464484
transform 1 0 37352 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_406
timestamp 1666464484
transform 1 0 38456 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_418
timestamp 1666464484
transform 1 0 39560 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_423
timestamp 1666464484
transform 1 0 40020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_435
timestamp 1666464484
transform 1 0 41124 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_447
timestamp 1666464484
transform 1 0 42228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_459
timestamp 1666464484
transform 1 0 43332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_471
timestamp 1666464484
transform 1 0 44436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_483
timestamp 1666464484
transform 1 0 45540 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_488
timestamp 1666464484
transform 1 0 46000 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_500
timestamp 1666464484
transform 1 0 47104 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_512
timestamp 1666464484
transform 1 0 48208 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_524
timestamp 1666464484
transform 1 0 49312 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_536
timestamp 1666464484
transform 1 0 50416 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_548
timestamp 1666464484
transform 1 0 51520 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_553
timestamp 1666464484
transform 1 0 51980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_565
timestamp 1666464484
transform 1 0 53084 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_577
timestamp 1666464484
transform 1 0 54188 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1666464484
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1666464484
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_613
timestamp 1666464484
transform 1 0 57500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_618
timestamp 1666464484
transform 1 0 57960 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_624
timestamp 1666464484
transform 1 0 58512 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1666464484
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1666464484
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_51
timestamp 1666464484
transform 1 0 5796 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_63
timestamp 1666464484
transform 1 0 6900 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_66
timestamp 1666464484
transform 1 0 7176 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_78
timestamp 1666464484
transform 1 0 8280 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_90
timestamp 1666464484
transform 1 0 9384 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_102
timestamp 1666464484
transform 1 0 10488 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_114
timestamp 1666464484
transform 1 0 11592 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_126
timestamp 1666464484
transform 1 0 12696 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_131
timestamp 1666464484
transform 1 0 13156 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_143
timestamp 1666464484
transform 1 0 14260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_155
timestamp 1666464484
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_179
timestamp 1666464484
transform 1 0 17572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_191
timestamp 1666464484
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_196
timestamp 1666464484
transform 1 0 19136 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_208
timestamp 1666464484
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_220
timestamp 1666464484
transform 1 0 21344 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_232
timestamp 1666464484
transform 1 0 22448 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_244
timestamp 1666464484
transform 1 0 23552 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_256
timestamp 1666464484
transform 1 0 24656 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666464484
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_285
timestamp 1666464484
transform 1 0 27324 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_297
timestamp 1666464484
transform 1 0 28428 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_309
timestamp 1666464484
transform 1 0 29532 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_321
timestamp 1666464484
transform 1 0 30636 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_326
timestamp 1666464484
transform 1 0 31096 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_338
timestamp 1666464484
transform 1 0 32200 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_350
timestamp 1666464484
transform 1 0 33304 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_362
timestamp 1666464484
transform 1 0 34408 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_374
timestamp 1666464484
transform 1 0 35512 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_386
timestamp 1666464484
transform 1 0 36616 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_391
timestamp 1666464484
transform 1 0 37076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_403
timestamp 1666464484
transform 1 0 38180 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_415
timestamp 1666464484
transform 1 0 39284 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_427
timestamp 1666464484
transform 1 0 40388 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_439
timestamp 1666464484
transform 1 0 41492 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_451
timestamp 1666464484
transform 1 0 42596 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_456
timestamp 1666464484
transform 1 0 43056 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_468
timestamp 1666464484
transform 1 0 44160 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_480
timestamp 1666464484
transform 1 0 45264 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_492
timestamp 1666464484
transform 1 0 46368 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_504
timestamp 1666464484
transform 1 0 47472 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_516
timestamp 1666464484
transform 1 0 48576 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_521
timestamp 1666464484
transform 1 0 49036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_533
timestamp 1666464484
transform 1 0 50140 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_545
timestamp 1666464484
transform 1 0 51244 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_557
timestamp 1666464484
transform 1 0 52348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_569
timestamp 1666464484
transform 1 0 53452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_581
timestamp 1666464484
transform 1 0 54556 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_586
timestamp 1666464484
transform 1 0 55016 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_598
timestamp 1666464484
transform 1 0 56120 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_610
timestamp 1666464484
transform 1 0 57224 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_622
timestamp 1666464484
transform 1 0 58328 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1666464484
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_31
timestamp 1666464484
transform 1 0 3956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_33
timestamp 1666464484
transform 1 0 4140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_45
timestamp 1666464484
transform 1 0 5244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_57
timestamp 1666464484
transform 1 0 6348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_69
timestamp 1666464484
transform 1 0 7452 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_81
timestamp 1666464484
transform 1 0 8556 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1666464484
transform 1 0 9660 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_98
timestamp 1666464484
transform 1 0 10120 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_110
timestamp 1666464484
transform 1 0 11224 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_122
timestamp 1666464484
transform 1 0 12328 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_134
timestamp 1666464484
transform 1 0 13432 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_146
timestamp 1666464484
transform 1 0 14536 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_158
timestamp 1666464484
transform 1 0 15640 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_163
timestamp 1666464484
transform 1 0 16100 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_175
timestamp 1666464484
transform 1 0 17204 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_187
timestamp 1666464484
transform 1 0 18308 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_199
timestamp 1666464484
transform 1 0 19412 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_211
timestamp 1666464484
transform 1 0 20516 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_223
timestamp 1666464484
transform 1 0 21620 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_228
timestamp 1666464484
transform 1 0 22080 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_240
timestamp 1666464484
transform 1 0 23184 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_252
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_264
timestamp 1666464484
transform 1 0 25392 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_276
timestamp 1666464484
transform 1 0 26496 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_288
timestamp 1666464484
transform 1 0 27600 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_293
timestamp 1666464484
transform 1 0 28060 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_305
timestamp 1666464484
transform 1 0 29164 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_317
timestamp 1666464484
transform 1 0 30268 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_329
timestamp 1666464484
transform 1 0 31372 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_341
timestamp 1666464484
transform 1 0 32476 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_353
timestamp 1666464484
transform 1 0 33580 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_358
timestamp 1666464484
transform 1 0 34040 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_370
timestamp 1666464484
transform 1 0 35144 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_382
timestamp 1666464484
transform 1 0 36248 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_394
timestamp 1666464484
transform 1 0 37352 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_406
timestamp 1666464484
transform 1 0 38456 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_418
timestamp 1666464484
transform 1 0 39560 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_423
timestamp 1666464484
transform 1 0 40020 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_435
timestamp 1666464484
transform 1 0 41124 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_447
timestamp 1666464484
transform 1 0 42228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_459
timestamp 1666464484
transform 1 0 43332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_471
timestamp 1666464484
transform 1 0 44436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_483
timestamp 1666464484
transform 1 0 45540 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_488
timestamp 1666464484
transform 1 0 46000 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_500
timestamp 1666464484
transform 1 0 47104 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_512
timestamp 1666464484
transform 1 0 48208 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_524
timestamp 1666464484
transform 1 0 49312 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_536
timestamp 1666464484
transform 1 0 50416 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_548
timestamp 1666464484
transform 1 0 51520 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_553
timestamp 1666464484
transform 1 0 51980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_565
timestamp 1666464484
transform 1 0 53084 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_577
timestamp 1666464484
transform 1 0 54188 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1666464484
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1666464484
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_613
timestamp 1666464484
transform 1 0 57500 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_618
timestamp 1666464484
transform 1 0 57960 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_624
timestamp 1666464484
transform 1 0 58512 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666464484
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_51
timestamp 1666464484
transform 1 0 5796 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_63
timestamp 1666464484
transform 1 0 6900 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_66
timestamp 1666464484
transform 1 0 7176 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_78
timestamp 1666464484
transform 1 0 8280 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_90
timestamp 1666464484
transform 1 0 9384 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_102
timestamp 1666464484
transform 1 0 10488 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_114
timestamp 1666464484
transform 1 0 11592 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_126
timestamp 1666464484
transform 1 0 12696 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_131
timestamp 1666464484
transform 1 0 13156 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_143
timestamp 1666464484
transform 1 0 14260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_155
timestamp 1666464484
transform 1 0 15364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_179
timestamp 1666464484
transform 1 0 17572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_191
timestamp 1666464484
transform 1 0 18676 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_196
timestamp 1666464484
transform 1 0 19136 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_208
timestamp 1666464484
transform 1 0 20240 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_220
timestamp 1666464484
transform 1 0 21344 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_232
timestamp 1666464484
transform 1 0 22448 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_244
timestamp 1666464484
transform 1 0 23552 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_256
timestamp 1666464484
transform 1 0 24656 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666464484
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_273
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_285
timestamp 1666464484
transform 1 0 27324 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_297
timestamp 1666464484
transform 1 0 28428 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_309
timestamp 1666464484
transform 1 0 29532 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_321
timestamp 1666464484
transform 1 0 30636 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_326
timestamp 1666464484
transform 1 0 31096 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_338
timestamp 1666464484
transform 1 0 32200 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_350
timestamp 1666464484
transform 1 0 33304 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_362
timestamp 1666464484
transform 1 0 34408 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_374
timestamp 1666464484
transform 1 0 35512 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_386
timestamp 1666464484
transform 1 0 36616 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_391
timestamp 1666464484
transform 1 0 37076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_403
timestamp 1666464484
transform 1 0 38180 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_415
timestamp 1666464484
transform 1 0 39284 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_427
timestamp 1666464484
transform 1 0 40388 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_439
timestamp 1666464484
transform 1 0 41492 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_451
timestamp 1666464484
transform 1 0 42596 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_456
timestamp 1666464484
transform 1 0 43056 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_468
timestamp 1666464484
transform 1 0 44160 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_480
timestamp 1666464484
transform 1 0 45264 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_492
timestamp 1666464484
transform 1 0 46368 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_504
timestamp 1666464484
transform 1 0 47472 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_516
timestamp 1666464484
transform 1 0 48576 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_521
timestamp 1666464484
transform 1 0 49036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_533
timestamp 1666464484
transform 1 0 50140 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_545
timestamp 1666464484
transform 1 0 51244 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_557
timestamp 1666464484
transform 1 0 52348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_569
timestamp 1666464484
transform 1 0 53452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_581
timestamp 1666464484
transform 1 0 54556 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_586
timestamp 1666464484
transform 1 0 55016 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_598
timestamp 1666464484
transform 1 0 56120 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_610
timestamp 1666464484
transform 1 0 57224 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_622
timestamp 1666464484
transform 1 0 58328 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_31
timestamp 1666464484
transform 1 0 3956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_33
timestamp 1666464484
transform 1 0 4140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_45
timestamp 1666464484
transform 1 0 5244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_57
timestamp 1666464484
transform 1 0 6348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_69
timestamp 1666464484
transform 1 0 7452 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_81
timestamp 1666464484
transform 1 0 8556 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1666464484
transform 1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_98
timestamp 1666464484
transform 1 0 10120 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_110
timestamp 1666464484
transform 1 0 11224 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_122
timestamp 1666464484
transform 1 0 12328 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_134
timestamp 1666464484
transform 1 0 13432 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_146
timestamp 1666464484
transform 1 0 14536 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_158
timestamp 1666464484
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_163
timestamp 1666464484
transform 1 0 16100 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_175
timestamp 1666464484
transform 1 0 17204 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_187
timestamp 1666464484
transform 1 0 18308 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_199
timestamp 1666464484
transform 1 0 19412 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_211
timestamp 1666464484
transform 1 0 20516 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_223
timestamp 1666464484
transform 1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_228
timestamp 1666464484
transform 1 0 22080 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_240
timestamp 1666464484
transform 1 0 23184 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_252
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_264
timestamp 1666464484
transform 1 0 25392 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_276
timestamp 1666464484
transform 1 0 26496 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_288
timestamp 1666464484
transform 1 0 27600 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_293
timestamp 1666464484
transform 1 0 28060 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_305
timestamp 1666464484
transform 1 0 29164 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_317
timestamp 1666464484
transform 1 0 30268 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_329
timestamp 1666464484
transform 1 0 31372 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_341
timestamp 1666464484
transform 1 0 32476 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_353
timestamp 1666464484
transform 1 0 33580 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_358
timestamp 1666464484
transform 1 0 34040 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_370
timestamp 1666464484
transform 1 0 35144 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_382
timestamp 1666464484
transform 1 0 36248 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_394
timestamp 1666464484
transform 1 0 37352 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_406
timestamp 1666464484
transform 1 0 38456 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_418
timestamp 1666464484
transform 1 0 39560 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_423
timestamp 1666464484
transform 1 0 40020 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_435
timestamp 1666464484
transform 1 0 41124 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_447
timestamp 1666464484
transform 1 0 42228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_459
timestamp 1666464484
transform 1 0 43332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_471
timestamp 1666464484
transform 1 0 44436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_483
timestamp 1666464484
transform 1 0 45540 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_488
timestamp 1666464484
transform 1 0 46000 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_500
timestamp 1666464484
transform 1 0 47104 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_512
timestamp 1666464484
transform 1 0 48208 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_524
timestamp 1666464484
transform 1 0 49312 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_536
timestamp 1666464484
transform 1 0 50416 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_548
timestamp 1666464484
transform 1 0 51520 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_553
timestamp 1666464484
transform 1 0 51980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_565
timestamp 1666464484
transform 1 0 53084 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_577
timestamp 1666464484
transform 1 0 54188 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1666464484
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1666464484
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_613
timestamp 1666464484
transform 1 0 57500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_618
timestamp 1666464484
transform 1 0 57960 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_624
timestamp 1666464484
transform 1 0 58512 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666464484
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1666464484
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_51
timestamp 1666464484
transform 1 0 5796 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_63
timestamp 1666464484
transform 1 0 6900 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_66
timestamp 1666464484
transform 1 0 7176 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_78
timestamp 1666464484
transform 1 0 8280 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_90
timestamp 1666464484
transform 1 0 9384 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_102
timestamp 1666464484
transform 1 0 10488 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_114
timestamp 1666464484
transform 1 0 11592 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_126
timestamp 1666464484
transform 1 0 12696 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_131
timestamp 1666464484
transform 1 0 13156 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_143
timestamp 1666464484
transform 1 0 14260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_155
timestamp 1666464484
transform 1 0 15364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_179
timestamp 1666464484
transform 1 0 17572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_191
timestamp 1666464484
transform 1 0 18676 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_196
timestamp 1666464484
transform 1 0 19136 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_208
timestamp 1666464484
transform 1 0 20240 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_220
timestamp 1666464484
transform 1 0 21344 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_232
timestamp 1666464484
transform 1 0 22448 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_244
timestamp 1666464484
transform 1 0 23552 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_256
timestamp 1666464484
transform 1 0 24656 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1666464484
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_273
timestamp 1666464484
transform 1 0 26220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_285
timestamp 1666464484
transform 1 0 27324 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_297
timestamp 1666464484
transform 1 0 28428 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_309
timestamp 1666464484
transform 1 0 29532 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_321
timestamp 1666464484
transform 1 0 30636 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_326
timestamp 1666464484
transform 1 0 31096 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_338
timestamp 1666464484
transform 1 0 32200 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_350
timestamp 1666464484
transform 1 0 33304 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_362
timestamp 1666464484
transform 1 0 34408 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_374
timestamp 1666464484
transform 1 0 35512 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_386
timestamp 1666464484
transform 1 0 36616 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_391
timestamp 1666464484
transform 1 0 37076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_403
timestamp 1666464484
transform 1 0 38180 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_415
timestamp 1666464484
transform 1 0 39284 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_427
timestamp 1666464484
transform 1 0 40388 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_439
timestamp 1666464484
transform 1 0 41492 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_451
timestamp 1666464484
transform 1 0 42596 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_456
timestamp 1666464484
transform 1 0 43056 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_468
timestamp 1666464484
transform 1 0 44160 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_480
timestamp 1666464484
transform 1 0 45264 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_492
timestamp 1666464484
transform 1 0 46368 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_504
timestamp 1666464484
transform 1 0 47472 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_516
timestamp 1666464484
transform 1 0 48576 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_521
timestamp 1666464484
transform 1 0 49036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_533
timestamp 1666464484
transform 1 0 50140 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_545
timestamp 1666464484
transform 1 0 51244 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_557
timestamp 1666464484
transform 1 0 52348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_569
timestamp 1666464484
transform 1 0 53452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_581
timestamp 1666464484
transform 1 0 54556 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_586
timestamp 1666464484
transform 1 0 55016 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_598
timestamp 1666464484
transform 1 0 56120 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_610
timestamp 1666464484
transform 1 0 57224 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_622
timestamp 1666464484
transform 1 0 58328 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_31
timestamp 1666464484
transform 1 0 3956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_33
timestamp 1666464484
transform 1 0 4140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_45
timestamp 1666464484
transform 1 0 5244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_57
timestamp 1666464484
transform 1 0 6348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_69
timestamp 1666464484
transform 1 0 7452 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_81
timestamp 1666464484
transform 1 0 8556 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1666464484
transform 1 0 9660 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_98
timestamp 1666464484
transform 1 0 10120 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_110
timestamp 1666464484
transform 1 0 11224 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_122
timestamp 1666464484
transform 1 0 12328 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_134
timestamp 1666464484
transform 1 0 13432 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_146
timestamp 1666464484
transform 1 0 14536 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_158
timestamp 1666464484
transform 1 0 15640 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_163
timestamp 1666464484
transform 1 0 16100 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_175
timestamp 1666464484
transform 1 0 17204 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_187
timestamp 1666464484
transform 1 0 18308 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_199
timestamp 1666464484
transform 1 0 19412 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_211
timestamp 1666464484
transform 1 0 20516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_223
timestamp 1666464484
transform 1 0 21620 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_228
timestamp 1666464484
transform 1 0 22080 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_240
timestamp 1666464484
transform 1 0 23184 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_252
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_264
timestamp 1666464484
transform 1 0 25392 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_276
timestamp 1666464484
transform 1 0 26496 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_288
timestamp 1666464484
transform 1 0 27600 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_293
timestamp 1666464484
transform 1 0 28060 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_305
timestamp 1666464484
transform 1 0 29164 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_317
timestamp 1666464484
transform 1 0 30268 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_329
timestamp 1666464484
transform 1 0 31372 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_341
timestamp 1666464484
transform 1 0 32476 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_353
timestamp 1666464484
transform 1 0 33580 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_358
timestamp 1666464484
transform 1 0 34040 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_370
timestamp 1666464484
transform 1 0 35144 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_382
timestamp 1666464484
transform 1 0 36248 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_394
timestamp 1666464484
transform 1 0 37352 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_406
timestamp 1666464484
transform 1 0 38456 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_418
timestamp 1666464484
transform 1 0 39560 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_423
timestamp 1666464484
transform 1 0 40020 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_435
timestamp 1666464484
transform 1 0 41124 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_447
timestamp 1666464484
transform 1 0 42228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_459
timestamp 1666464484
transform 1 0 43332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_471
timestamp 1666464484
transform 1 0 44436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_483
timestamp 1666464484
transform 1 0 45540 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_488
timestamp 1666464484
transform 1 0 46000 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_500
timestamp 1666464484
transform 1 0 47104 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_512
timestamp 1666464484
transform 1 0 48208 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_524
timestamp 1666464484
transform 1 0 49312 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_536
timestamp 1666464484
transform 1 0 50416 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_548
timestamp 1666464484
transform 1 0 51520 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_553
timestamp 1666464484
transform 1 0 51980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_565
timestamp 1666464484
transform 1 0 53084 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_577
timestamp 1666464484
transform 1 0 54188 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1666464484
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1666464484
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_613
timestamp 1666464484
transform 1 0 57500 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_618
timestamp 1666464484
transform 1 0 57960 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_624
timestamp 1666464484
transform 1 0 58512 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_51
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_63
timestamp 1666464484
transform 1 0 6900 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_66
timestamp 1666464484
transform 1 0 7176 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_78
timestamp 1666464484
transform 1 0 8280 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_90
timestamp 1666464484
transform 1 0 9384 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_102
timestamp 1666464484
transform 1 0 10488 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_114
timestamp 1666464484
transform 1 0 11592 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_126
timestamp 1666464484
transform 1 0 12696 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_131
timestamp 1666464484
transform 1 0 13156 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_143
timestamp 1666464484
transform 1 0 14260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_155
timestamp 1666464484
transform 1 0 15364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_179
timestamp 1666464484
transform 1 0 17572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_191
timestamp 1666464484
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_196
timestamp 1666464484
transform 1 0 19136 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_208
timestamp 1666464484
transform 1 0 20240 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_220
timestamp 1666464484
transform 1 0 21344 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_232
timestamp 1666464484
transform 1 0 22448 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_244
timestamp 1666464484
transform 1 0 23552 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_256
timestamp 1666464484
transform 1 0 24656 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666464484
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_273
timestamp 1666464484
transform 1 0 26220 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_285
timestamp 1666464484
transform 1 0 27324 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_297
timestamp 1666464484
transform 1 0 28428 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_309
timestamp 1666464484
transform 1 0 29532 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_321
timestamp 1666464484
transform 1 0 30636 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_326
timestamp 1666464484
transform 1 0 31096 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_338
timestamp 1666464484
transform 1 0 32200 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_350
timestamp 1666464484
transform 1 0 33304 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_362
timestamp 1666464484
transform 1 0 34408 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_374
timestamp 1666464484
transform 1 0 35512 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_386
timestamp 1666464484
transform 1 0 36616 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_391
timestamp 1666464484
transform 1 0 37076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_403
timestamp 1666464484
transform 1 0 38180 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_415
timestamp 1666464484
transform 1 0 39284 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_427
timestamp 1666464484
transform 1 0 40388 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_439
timestamp 1666464484
transform 1 0 41492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_451
timestamp 1666464484
transform 1 0 42596 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_456
timestamp 1666464484
transform 1 0 43056 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_468
timestamp 1666464484
transform 1 0 44160 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_480
timestamp 1666464484
transform 1 0 45264 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_492
timestamp 1666464484
transform 1 0 46368 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_504
timestamp 1666464484
transform 1 0 47472 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_516
timestamp 1666464484
transform 1 0 48576 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_521
timestamp 1666464484
transform 1 0 49036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_533
timestamp 1666464484
transform 1 0 50140 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_545
timestamp 1666464484
transform 1 0 51244 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_557
timestamp 1666464484
transform 1 0 52348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_569
timestamp 1666464484
transform 1 0 53452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_581
timestamp 1666464484
transform 1 0 54556 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_586
timestamp 1666464484
transform 1 0 55016 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_598
timestamp 1666464484
transform 1 0 56120 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_610
timestamp 1666464484
transform 1 0 57224 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_622
timestamp 1666464484
transform 1 0 58328 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1666464484
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1666464484
transform 1 0 3588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_31
timestamp 1666464484
transform 1 0 3956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_33
timestamp 1666464484
transform 1 0 4140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_45
timestamp 1666464484
transform 1 0 5244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_57
timestamp 1666464484
transform 1 0 6348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_69
timestamp 1666464484
transform 1 0 7452 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_81
timestamp 1666464484
transform 1 0 8556 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_93
timestamp 1666464484
transform 1 0 9660 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_98
timestamp 1666464484
transform 1 0 10120 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_110
timestamp 1666464484
transform 1 0 11224 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_122
timestamp 1666464484
transform 1 0 12328 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_134
timestamp 1666464484
transform 1 0 13432 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_146
timestamp 1666464484
transform 1 0 14536 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_158
timestamp 1666464484
transform 1 0 15640 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_163
timestamp 1666464484
transform 1 0 16100 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_175
timestamp 1666464484
transform 1 0 17204 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_187
timestamp 1666464484
transform 1 0 18308 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_199
timestamp 1666464484
transform 1 0 19412 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_211
timestamp 1666464484
transform 1 0 20516 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_223
timestamp 1666464484
transform 1 0 21620 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_228
timestamp 1666464484
transform 1 0 22080 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_240
timestamp 1666464484
transform 1 0 23184 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_252
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_264
timestamp 1666464484
transform 1 0 25392 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_276
timestamp 1666464484
transform 1 0 26496 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_288
timestamp 1666464484
transform 1 0 27600 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_293
timestamp 1666464484
transform 1 0 28060 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_305
timestamp 1666464484
transform 1 0 29164 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_317
timestamp 1666464484
transform 1 0 30268 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_329
timestamp 1666464484
transform 1 0 31372 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_341
timestamp 1666464484
transform 1 0 32476 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_353
timestamp 1666464484
transform 1 0 33580 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_358
timestamp 1666464484
transform 1 0 34040 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_370
timestamp 1666464484
transform 1 0 35144 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_382
timestamp 1666464484
transform 1 0 36248 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_394
timestamp 1666464484
transform 1 0 37352 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_406
timestamp 1666464484
transform 1 0 38456 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_418
timestamp 1666464484
transform 1 0 39560 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_423
timestamp 1666464484
transform 1 0 40020 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_435
timestamp 1666464484
transform 1 0 41124 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_447
timestamp 1666464484
transform 1 0 42228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_459
timestamp 1666464484
transform 1 0 43332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_471
timestamp 1666464484
transform 1 0 44436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_483
timestamp 1666464484
transform 1 0 45540 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_488
timestamp 1666464484
transform 1 0 46000 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_500
timestamp 1666464484
transform 1 0 47104 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_512
timestamp 1666464484
transform 1 0 48208 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_524
timestamp 1666464484
transform 1 0 49312 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_536
timestamp 1666464484
transform 1 0 50416 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_548
timestamp 1666464484
transform 1 0 51520 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_553
timestamp 1666464484
transform 1 0 51980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_565
timestamp 1666464484
transform 1 0 53084 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_577
timestamp 1666464484
transform 1 0 54188 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1666464484
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1666464484
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_613
timestamp 1666464484
transform 1 0 57500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_618
timestamp 1666464484
transform 1 0 57960 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_624
timestamp 1666464484
transform 1 0 58512 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_63
timestamp 1666464484
transform 1 0 6900 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_66
timestamp 1666464484
transform 1 0 7176 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_78
timestamp 1666464484
transform 1 0 8280 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_90
timestamp 1666464484
transform 1 0 9384 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_102
timestamp 1666464484
transform 1 0 10488 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_114
timestamp 1666464484
transform 1 0 11592 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_126
timestamp 1666464484
transform 1 0 12696 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_131
timestamp 1666464484
transform 1 0 13156 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_143
timestamp 1666464484
transform 1 0 14260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_155
timestamp 1666464484
transform 1 0 15364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_179
timestamp 1666464484
transform 1 0 17572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_191
timestamp 1666464484
transform 1 0 18676 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_196
timestamp 1666464484
transform 1 0 19136 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_208
timestamp 1666464484
transform 1 0 20240 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_220
timestamp 1666464484
transform 1 0 21344 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_232
timestamp 1666464484
transform 1 0 22448 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_244
timestamp 1666464484
transform 1 0 23552 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1666464484
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666464484
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_273
timestamp 1666464484
transform 1 0 26220 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_285
timestamp 1666464484
transform 1 0 27324 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_297
timestamp 1666464484
transform 1 0 28428 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_309
timestamp 1666464484
transform 1 0 29532 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_321
timestamp 1666464484
transform 1 0 30636 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_326
timestamp 1666464484
transform 1 0 31096 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_338
timestamp 1666464484
transform 1 0 32200 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_350
timestamp 1666464484
transform 1 0 33304 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_362
timestamp 1666464484
transform 1 0 34408 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_374
timestamp 1666464484
transform 1 0 35512 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_386
timestamp 1666464484
transform 1 0 36616 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_391
timestamp 1666464484
transform 1 0 37076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_403
timestamp 1666464484
transform 1 0 38180 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_415
timestamp 1666464484
transform 1 0 39284 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_427
timestamp 1666464484
transform 1 0 40388 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_439
timestamp 1666464484
transform 1 0 41492 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_451
timestamp 1666464484
transform 1 0 42596 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_456
timestamp 1666464484
transform 1 0 43056 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_468
timestamp 1666464484
transform 1 0 44160 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_480
timestamp 1666464484
transform 1 0 45264 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_492
timestamp 1666464484
transform 1 0 46368 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_504
timestamp 1666464484
transform 1 0 47472 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_516
timestamp 1666464484
transform 1 0 48576 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_521
timestamp 1666464484
transform 1 0 49036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_533
timestamp 1666464484
transform 1 0 50140 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_545
timestamp 1666464484
transform 1 0 51244 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_557
timestamp 1666464484
transform 1 0 52348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_569
timestamp 1666464484
transform 1 0 53452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_581
timestamp 1666464484
transform 1 0 54556 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_586
timestamp 1666464484
transform 1 0 55016 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_598
timestamp 1666464484
transform 1 0 56120 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_610
timestamp 1666464484
transform 1 0 57224 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_622
timestamp 1666464484
transform 1 0 58328 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1666464484
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_31
timestamp 1666464484
transform 1 0 3956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_33
timestamp 1666464484
transform 1 0 4140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_45
timestamp 1666464484
transform 1 0 5244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_57
timestamp 1666464484
transform 1 0 6348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_69
timestamp 1666464484
transform 1 0 7452 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_81
timestamp 1666464484
transform 1 0 8556 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_93
timestamp 1666464484
transform 1 0 9660 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_98
timestamp 1666464484
transform 1 0 10120 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_110
timestamp 1666464484
transform 1 0 11224 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_122
timestamp 1666464484
transform 1 0 12328 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_134
timestamp 1666464484
transform 1 0 13432 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_146
timestamp 1666464484
transform 1 0 14536 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_158
timestamp 1666464484
transform 1 0 15640 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_163
timestamp 1666464484
transform 1 0 16100 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_175
timestamp 1666464484
transform 1 0 17204 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_187
timestamp 1666464484
transform 1 0 18308 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_199
timestamp 1666464484
transform 1 0 19412 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_211
timestamp 1666464484
transform 1 0 20516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_223
timestamp 1666464484
transform 1 0 21620 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_228
timestamp 1666464484
transform 1 0 22080 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_240
timestamp 1666464484
transform 1 0 23184 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_252
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_264
timestamp 1666464484
transform 1 0 25392 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_276
timestamp 1666464484
transform 1 0 26496 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_288
timestamp 1666464484
transform 1 0 27600 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_293
timestamp 1666464484
transform 1 0 28060 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_305
timestamp 1666464484
transform 1 0 29164 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_317
timestamp 1666464484
transform 1 0 30268 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_329
timestamp 1666464484
transform 1 0 31372 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_341
timestamp 1666464484
transform 1 0 32476 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_353
timestamp 1666464484
transform 1 0 33580 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_358
timestamp 1666464484
transform 1 0 34040 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_370
timestamp 1666464484
transform 1 0 35144 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_382
timestamp 1666464484
transform 1 0 36248 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_394
timestamp 1666464484
transform 1 0 37352 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_406
timestamp 1666464484
transform 1 0 38456 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_418
timestamp 1666464484
transform 1 0 39560 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_423
timestamp 1666464484
transform 1 0 40020 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_435
timestamp 1666464484
transform 1 0 41124 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_447
timestamp 1666464484
transform 1 0 42228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_459
timestamp 1666464484
transform 1 0 43332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_471
timestamp 1666464484
transform 1 0 44436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_483
timestamp 1666464484
transform 1 0 45540 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_488
timestamp 1666464484
transform 1 0 46000 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_500
timestamp 1666464484
transform 1 0 47104 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_512
timestamp 1666464484
transform 1 0 48208 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_524
timestamp 1666464484
transform 1 0 49312 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_536
timestamp 1666464484
transform 1 0 50416 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_548
timestamp 1666464484
transform 1 0 51520 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_553
timestamp 1666464484
transform 1 0 51980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_565
timestamp 1666464484
transform 1 0 53084 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_577
timestamp 1666464484
transform 1 0 54188 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1666464484
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1666464484
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_613
timestamp 1666464484
transform 1 0 57500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_618
timestamp 1666464484
transform 1 0 57960 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_624
timestamp 1666464484
transform 1 0 58512 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666464484
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_51
timestamp 1666464484
transform 1 0 5796 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_63
timestamp 1666464484
transform 1 0 6900 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_66
timestamp 1666464484
transform 1 0 7176 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_78
timestamp 1666464484
transform 1 0 8280 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_90
timestamp 1666464484
transform 1 0 9384 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_102
timestamp 1666464484
transform 1 0 10488 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_114
timestamp 1666464484
transform 1 0 11592 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_126
timestamp 1666464484
transform 1 0 12696 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_131
timestamp 1666464484
transform 1 0 13156 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_143
timestamp 1666464484
transform 1 0 14260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_155
timestamp 1666464484
transform 1 0 15364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_179
timestamp 1666464484
transform 1 0 17572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_191
timestamp 1666464484
transform 1 0 18676 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_196
timestamp 1666464484
transform 1 0 19136 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_208
timestamp 1666464484
transform 1 0 20240 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_220
timestamp 1666464484
transform 1 0 21344 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_232
timestamp 1666464484
transform 1 0 22448 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_244
timestamp 1666464484
transform 1 0 23552 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_256
timestamp 1666464484
transform 1 0 24656 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1666464484
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_273
timestamp 1666464484
transform 1 0 26220 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_285
timestamp 1666464484
transform 1 0 27324 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_297
timestamp 1666464484
transform 1 0 28428 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_309
timestamp 1666464484
transform 1 0 29532 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_321
timestamp 1666464484
transform 1 0 30636 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_326
timestamp 1666464484
transform 1 0 31096 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_338
timestamp 1666464484
transform 1 0 32200 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_350
timestamp 1666464484
transform 1 0 33304 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_362
timestamp 1666464484
transform 1 0 34408 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_374
timestamp 1666464484
transform 1 0 35512 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_386
timestamp 1666464484
transform 1 0 36616 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_391
timestamp 1666464484
transform 1 0 37076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_403
timestamp 1666464484
transform 1 0 38180 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_415
timestamp 1666464484
transform 1 0 39284 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_427
timestamp 1666464484
transform 1 0 40388 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_439
timestamp 1666464484
transform 1 0 41492 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_451
timestamp 1666464484
transform 1 0 42596 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_456
timestamp 1666464484
transform 1 0 43056 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_468
timestamp 1666464484
transform 1 0 44160 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_480
timestamp 1666464484
transform 1 0 45264 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_492
timestamp 1666464484
transform 1 0 46368 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_504
timestamp 1666464484
transform 1 0 47472 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_516
timestamp 1666464484
transform 1 0 48576 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_521
timestamp 1666464484
transform 1 0 49036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_533
timestamp 1666464484
transform 1 0 50140 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_545
timestamp 1666464484
transform 1 0 51244 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_557
timestamp 1666464484
transform 1 0 52348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_569
timestamp 1666464484
transform 1 0 53452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_581
timestamp 1666464484
transform 1 0 54556 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_586
timestamp 1666464484
transform 1 0 55016 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_598
timestamp 1666464484
transform 1 0 56120 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_610
timestamp 1666464484
transform 1 0 57224 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_622
timestamp 1666464484
transform 1 0 58328 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_31
timestamp 1666464484
transform 1 0 3956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_33
timestamp 1666464484
transform 1 0 4140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_45
timestamp 1666464484
transform 1 0 5244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_57
timestamp 1666464484
transform 1 0 6348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_69
timestamp 1666464484
transform 1 0 7452 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_81
timestamp 1666464484
transform 1 0 8556 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1666464484
transform 1 0 9660 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_98
timestamp 1666464484
transform 1 0 10120 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_110
timestamp 1666464484
transform 1 0 11224 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_122
timestamp 1666464484
transform 1 0 12328 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_134
timestamp 1666464484
transform 1 0 13432 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_146
timestamp 1666464484
transform 1 0 14536 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_158
timestamp 1666464484
transform 1 0 15640 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_163
timestamp 1666464484
transform 1 0 16100 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_175
timestamp 1666464484
transform 1 0 17204 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_187
timestamp 1666464484
transform 1 0 18308 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_199
timestamp 1666464484
transform 1 0 19412 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_211
timestamp 1666464484
transform 1 0 20516 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_223
timestamp 1666464484
transform 1 0 21620 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_228
timestamp 1666464484
transform 1 0 22080 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_240
timestamp 1666464484
transform 1 0 23184 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_252
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_264
timestamp 1666464484
transform 1 0 25392 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_276
timestamp 1666464484
transform 1 0 26496 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_288
timestamp 1666464484
transform 1 0 27600 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_293
timestamp 1666464484
transform 1 0 28060 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_305
timestamp 1666464484
transform 1 0 29164 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_317
timestamp 1666464484
transform 1 0 30268 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_329
timestamp 1666464484
transform 1 0 31372 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_341
timestamp 1666464484
transform 1 0 32476 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_353
timestamp 1666464484
transform 1 0 33580 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_358
timestamp 1666464484
transform 1 0 34040 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_370
timestamp 1666464484
transform 1 0 35144 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_382
timestamp 1666464484
transform 1 0 36248 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_394
timestamp 1666464484
transform 1 0 37352 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_406
timestamp 1666464484
transform 1 0 38456 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_418
timestamp 1666464484
transform 1 0 39560 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_423
timestamp 1666464484
transform 1 0 40020 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_435
timestamp 1666464484
transform 1 0 41124 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_447
timestamp 1666464484
transform 1 0 42228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_459
timestamp 1666464484
transform 1 0 43332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_471
timestamp 1666464484
transform 1 0 44436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_483
timestamp 1666464484
transform 1 0 45540 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_488
timestamp 1666464484
transform 1 0 46000 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_500
timestamp 1666464484
transform 1 0 47104 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_512
timestamp 1666464484
transform 1 0 48208 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_524
timestamp 1666464484
transform 1 0 49312 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_536
timestamp 1666464484
transform 1 0 50416 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_548
timestamp 1666464484
transform 1 0 51520 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_553
timestamp 1666464484
transform 1 0 51980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_565
timestamp 1666464484
transform 1 0 53084 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_577
timestamp 1666464484
transform 1 0 54188 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1666464484
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1666464484
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_613
timestamp 1666464484
transform 1 0 57500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_618
timestamp 1666464484
transform 1 0 57960 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_624
timestamp 1666464484
transform 1 0 58512 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1666464484
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_51
timestamp 1666464484
transform 1 0 5796 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_63
timestamp 1666464484
transform 1 0 6900 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_66
timestamp 1666464484
transform 1 0 7176 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_78
timestamp 1666464484
transform 1 0 8280 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_90
timestamp 1666464484
transform 1 0 9384 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_102
timestamp 1666464484
transform 1 0 10488 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_114
timestamp 1666464484
transform 1 0 11592 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_126
timestamp 1666464484
transform 1 0 12696 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_131
timestamp 1666464484
transform 1 0 13156 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_143
timestamp 1666464484
transform 1 0 14260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_155
timestamp 1666464484
transform 1 0 15364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_179
timestamp 1666464484
transform 1 0 17572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_191
timestamp 1666464484
transform 1 0 18676 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_196
timestamp 1666464484
transform 1 0 19136 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_208
timestamp 1666464484
transform 1 0 20240 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_220
timestamp 1666464484
transform 1 0 21344 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_232
timestamp 1666464484
transform 1 0 22448 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_244
timestamp 1666464484
transform 1 0 23552 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_256
timestamp 1666464484
transform 1 0 24656 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1666464484
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_273
timestamp 1666464484
transform 1 0 26220 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_285
timestamp 1666464484
transform 1 0 27324 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_297
timestamp 1666464484
transform 1 0 28428 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_309
timestamp 1666464484
transform 1 0 29532 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_321
timestamp 1666464484
transform 1 0 30636 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_326
timestamp 1666464484
transform 1 0 31096 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_338
timestamp 1666464484
transform 1 0 32200 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_350
timestamp 1666464484
transform 1 0 33304 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_362
timestamp 1666464484
transform 1 0 34408 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_374
timestamp 1666464484
transform 1 0 35512 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_386
timestamp 1666464484
transform 1 0 36616 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_391
timestamp 1666464484
transform 1 0 37076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_403
timestamp 1666464484
transform 1 0 38180 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_415
timestamp 1666464484
transform 1 0 39284 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_427
timestamp 1666464484
transform 1 0 40388 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_439
timestamp 1666464484
transform 1 0 41492 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_451
timestamp 1666464484
transform 1 0 42596 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_456
timestamp 1666464484
transform 1 0 43056 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_468
timestamp 1666464484
transform 1 0 44160 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_480
timestamp 1666464484
transform 1 0 45264 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_492
timestamp 1666464484
transform 1 0 46368 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_504
timestamp 1666464484
transform 1 0 47472 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_516
timestamp 1666464484
transform 1 0 48576 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_521
timestamp 1666464484
transform 1 0 49036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_533
timestamp 1666464484
transform 1 0 50140 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_545
timestamp 1666464484
transform 1 0 51244 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_557
timestamp 1666464484
transform 1 0 52348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_569
timestamp 1666464484
transform 1 0 53452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_581
timestamp 1666464484
transform 1 0 54556 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_586
timestamp 1666464484
transform 1 0 55016 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_598
timestamp 1666464484
transform 1 0 56120 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_610
timestamp 1666464484
transform 1 0 57224 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_622
timestamp 1666464484
transform 1 0 58328 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_31
timestamp 1666464484
transform 1 0 3956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_33
timestamp 1666464484
transform 1 0 4140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_45
timestamp 1666464484
transform 1 0 5244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_57
timestamp 1666464484
transform 1 0 6348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_69
timestamp 1666464484
transform 1 0 7452 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_81
timestamp 1666464484
transform 1 0 8556 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1666464484
transform 1 0 9660 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_98
timestamp 1666464484
transform 1 0 10120 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_110
timestamp 1666464484
transform 1 0 11224 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_122
timestamp 1666464484
transform 1 0 12328 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_134
timestamp 1666464484
transform 1 0 13432 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_146
timestamp 1666464484
transform 1 0 14536 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_158
timestamp 1666464484
transform 1 0 15640 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_163
timestamp 1666464484
transform 1 0 16100 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_175
timestamp 1666464484
transform 1 0 17204 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_187
timestamp 1666464484
transform 1 0 18308 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_199
timestamp 1666464484
transform 1 0 19412 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_211
timestamp 1666464484
transform 1 0 20516 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_223
timestamp 1666464484
transform 1 0 21620 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_228
timestamp 1666464484
transform 1 0 22080 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_240
timestamp 1666464484
transform 1 0 23184 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_252
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_264
timestamp 1666464484
transform 1 0 25392 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_276
timestamp 1666464484
transform 1 0 26496 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_288
timestamp 1666464484
transform 1 0 27600 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_293
timestamp 1666464484
transform 1 0 28060 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_305
timestamp 1666464484
transform 1 0 29164 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_317
timestamp 1666464484
transform 1 0 30268 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_329
timestamp 1666464484
transform 1 0 31372 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_341
timestamp 1666464484
transform 1 0 32476 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_353
timestamp 1666464484
transform 1 0 33580 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_358
timestamp 1666464484
transform 1 0 34040 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_370
timestamp 1666464484
transform 1 0 35144 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_382
timestamp 1666464484
transform 1 0 36248 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_394
timestamp 1666464484
transform 1 0 37352 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_406
timestamp 1666464484
transform 1 0 38456 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_418
timestamp 1666464484
transform 1 0 39560 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_423
timestamp 1666464484
transform 1 0 40020 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_435
timestamp 1666464484
transform 1 0 41124 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_447
timestamp 1666464484
transform 1 0 42228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_459
timestamp 1666464484
transform 1 0 43332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_471
timestamp 1666464484
transform 1 0 44436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_483
timestamp 1666464484
transform 1 0 45540 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_488
timestamp 1666464484
transform 1 0 46000 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_500
timestamp 1666464484
transform 1 0 47104 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_512
timestamp 1666464484
transform 1 0 48208 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_524
timestamp 1666464484
transform 1 0 49312 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_536
timestamp 1666464484
transform 1 0 50416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_548
timestamp 1666464484
transform 1 0 51520 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_553
timestamp 1666464484
transform 1 0 51980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_565
timestamp 1666464484
transform 1 0 53084 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_577
timestamp 1666464484
transform 1 0 54188 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1666464484
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1666464484
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_613
timestamp 1666464484
transform 1 0 57500 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_618
timestamp 1666464484
transform 1 0 57960 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_624
timestamp 1666464484
transform 1 0 58512 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_51
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_63
timestamp 1666464484
transform 1 0 6900 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_66
timestamp 1666464484
transform 1 0 7176 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_78
timestamp 1666464484
transform 1 0 8280 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_90
timestamp 1666464484
transform 1 0 9384 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_102
timestamp 1666464484
transform 1 0 10488 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_114
timestamp 1666464484
transform 1 0 11592 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_126
timestamp 1666464484
transform 1 0 12696 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_131
timestamp 1666464484
transform 1 0 13156 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_143
timestamp 1666464484
transform 1 0 14260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_155
timestamp 1666464484
transform 1 0 15364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_179
timestamp 1666464484
transform 1 0 17572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_191
timestamp 1666464484
transform 1 0 18676 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_196
timestamp 1666464484
transform 1 0 19136 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_208
timestamp 1666464484
transform 1 0 20240 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_220
timestamp 1666464484
transform 1 0 21344 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_232
timestamp 1666464484
transform 1 0 22448 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_244
timestamp 1666464484
transform 1 0 23552 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_256
timestamp 1666464484
transform 1 0 24656 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1666464484
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_273
timestamp 1666464484
transform 1 0 26220 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_285
timestamp 1666464484
transform 1 0 27324 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_297
timestamp 1666464484
transform 1 0 28428 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_309
timestamp 1666464484
transform 1 0 29532 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_321
timestamp 1666464484
transform 1 0 30636 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_326
timestamp 1666464484
transform 1 0 31096 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_338
timestamp 1666464484
transform 1 0 32200 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_350
timestamp 1666464484
transform 1 0 33304 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_362
timestamp 1666464484
transform 1 0 34408 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_374
timestamp 1666464484
transform 1 0 35512 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_386
timestamp 1666464484
transform 1 0 36616 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_391
timestamp 1666464484
transform 1 0 37076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_403
timestamp 1666464484
transform 1 0 38180 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_415
timestamp 1666464484
transform 1 0 39284 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_427
timestamp 1666464484
transform 1 0 40388 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_439
timestamp 1666464484
transform 1 0 41492 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_451
timestamp 1666464484
transform 1 0 42596 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_456
timestamp 1666464484
transform 1 0 43056 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_468
timestamp 1666464484
transform 1 0 44160 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_480
timestamp 1666464484
transform 1 0 45264 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_492
timestamp 1666464484
transform 1 0 46368 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_504
timestamp 1666464484
transform 1 0 47472 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_516
timestamp 1666464484
transform 1 0 48576 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_521
timestamp 1666464484
transform 1 0 49036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_533
timestamp 1666464484
transform 1 0 50140 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_545
timestamp 1666464484
transform 1 0 51244 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_557
timestamp 1666464484
transform 1 0 52348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_569
timestamp 1666464484
transform 1 0 53452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_581
timestamp 1666464484
transform 1 0 54556 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_586
timestamp 1666464484
transform 1 0 55016 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_598
timestamp 1666464484
transform 1 0 56120 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_610
timestamp 1666464484
transform 1 0 57224 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_622
timestamp 1666464484
transform 1 0 58328 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1666464484
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1666464484
transform 1 0 3588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_31
timestamp 1666464484
transform 1 0 3956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_33
timestamp 1666464484
transform 1 0 4140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_45
timestamp 1666464484
transform 1 0 5244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_57
timestamp 1666464484
transform 1 0 6348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_69
timestamp 1666464484
transform 1 0 7452 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_81
timestamp 1666464484
transform 1 0 8556 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_93
timestamp 1666464484
transform 1 0 9660 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_98
timestamp 1666464484
transform 1 0 10120 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_110
timestamp 1666464484
transform 1 0 11224 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_122
timestamp 1666464484
transform 1 0 12328 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_134
timestamp 1666464484
transform 1 0 13432 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_146
timestamp 1666464484
transform 1 0 14536 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_158
timestamp 1666464484
transform 1 0 15640 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_163
timestamp 1666464484
transform 1 0 16100 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_175
timestamp 1666464484
transform 1 0 17204 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_187
timestamp 1666464484
transform 1 0 18308 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_199
timestamp 1666464484
transform 1 0 19412 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_211
timestamp 1666464484
transform 1 0 20516 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_223
timestamp 1666464484
transform 1 0 21620 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_228
timestamp 1666464484
transform 1 0 22080 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_240
timestamp 1666464484
transform 1 0 23184 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_252
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_264
timestamp 1666464484
transform 1 0 25392 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_276
timestamp 1666464484
transform 1 0 26496 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_288
timestamp 1666464484
transform 1 0 27600 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_293
timestamp 1666464484
transform 1 0 28060 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_305
timestamp 1666464484
transform 1 0 29164 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_317
timestamp 1666464484
transform 1 0 30268 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_329
timestamp 1666464484
transform 1 0 31372 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_341
timestamp 1666464484
transform 1 0 32476 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_353
timestamp 1666464484
transform 1 0 33580 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_358
timestamp 1666464484
transform 1 0 34040 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_370
timestamp 1666464484
transform 1 0 35144 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_382
timestamp 1666464484
transform 1 0 36248 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_394
timestamp 1666464484
transform 1 0 37352 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_406
timestamp 1666464484
transform 1 0 38456 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_418
timestamp 1666464484
transform 1 0 39560 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_423
timestamp 1666464484
transform 1 0 40020 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_435
timestamp 1666464484
transform 1 0 41124 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_447
timestamp 1666464484
transform 1 0 42228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_459
timestamp 1666464484
transform 1 0 43332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_471
timestamp 1666464484
transform 1 0 44436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_483
timestamp 1666464484
transform 1 0 45540 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_488
timestamp 1666464484
transform 1 0 46000 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_500
timestamp 1666464484
transform 1 0 47104 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_512
timestamp 1666464484
transform 1 0 48208 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_524
timestamp 1666464484
transform 1 0 49312 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_536
timestamp 1666464484
transform 1 0 50416 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_548
timestamp 1666464484
transform 1 0 51520 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_553
timestamp 1666464484
transform 1 0 51980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_565
timestamp 1666464484
transform 1 0 53084 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_577
timestamp 1666464484
transform 1 0 54188 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1666464484
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1666464484
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_613
timestamp 1666464484
transform 1 0 57500 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_618
timestamp 1666464484
transform 1 0 57960 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_624
timestamp 1666464484
transform 1 0 58512 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666464484
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1666464484
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1666464484
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_51
timestamp 1666464484
transform 1 0 5796 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_63
timestamp 1666464484
transform 1 0 6900 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_66
timestamp 1666464484
transform 1 0 7176 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_78
timestamp 1666464484
transform 1 0 8280 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_90
timestamp 1666464484
transform 1 0 9384 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_102
timestamp 1666464484
transform 1 0 10488 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_114
timestamp 1666464484
transform 1 0 11592 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_126
timestamp 1666464484
transform 1 0 12696 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_131
timestamp 1666464484
transform 1 0 13156 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_143
timestamp 1666464484
transform 1 0 14260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_155
timestamp 1666464484
transform 1 0 15364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_179
timestamp 1666464484
transform 1 0 17572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_191
timestamp 1666464484
transform 1 0 18676 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_196
timestamp 1666464484
transform 1 0 19136 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_208
timestamp 1666464484
transform 1 0 20240 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_220
timestamp 1666464484
transform 1 0 21344 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_232
timestamp 1666464484
transform 1 0 22448 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_244
timestamp 1666464484
transform 1 0 23552 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_256
timestamp 1666464484
transform 1 0 24656 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1666464484
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_273
timestamp 1666464484
transform 1 0 26220 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_285
timestamp 1666464484
transform 1 0 27324 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_297
timestamp 1666464484
transform 1 0 28428 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_309
timestamp 1666464484
transform 1 0 29532 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_321
timestamp 1666464484
transform 1 0 30636 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_326
timestamp 1666464484
transform 1 0 31096 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_338
timestamp 1666464484
transform 1 0 32200 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_350
timestamp 1666464484
transform 1 0 33304 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_362
timestamp 1666464484
transform 1 0 34408 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_374
timestamp 1666464484
transform 1 0 35512 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_386
timestamp 1666464484
transform 1 0 36616 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_391
timestamp 1666464484
transform 1 0 37076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_403
timestamp 1666464484
transform 1 0 38180 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_415
timestamp 1666464484
transform 1 0 39284 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_427
timestamp 1666464484
transform 1 0 40388 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_439
timestamp 1666464484
transform 1 0 41492 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_451
timestamp 1666464484
transform 1 0 42596 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_456
timestamp 1666464484
transform 1 0 43056 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_468
timestamp 1666464484
transform 1 0 44160 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_480
timestamp 1666464484
transform 1 0 45264 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_492
timestamp 1666464484
transform 1 0 46368 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_504
timestamp 1666464484
transform 1 0 47472 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_516
timestamp 1666464484
transform 1 0 48576 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_521
timestamp 1666464484
transform 1 0 49036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_533
timestamp 1666464484
transform 1 0 50140 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_545
timestamp 1666464484
transform 1 0 51244 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_557
timestamp 1666464484
transform 1 0 52348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_569
timestamp 1666464484
transform 1 0 53452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_581
timestamp 1666464484
transform 1 0 54556 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_586
timestamp 1666464484
transform 1 0 55016 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_598
timestamp 1666464484
transform 1 0 56120 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_610
timestamp 1666464484
transform 1 0 57224 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_622
timestamp 1666464484
transform 1 0 58328 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_31
timestamp 1666464484
transform 1 0 3956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_33
timestamp 1666464484
transform 1 0 4140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_45
timestamp 1666464484
transform 1 0 5244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_57
timestamp 1666464484
transform 1 0 6348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_69
timestamp 1666464484
transform 1 0 7452 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_81
timestamp 1666464484
transform 1 0 8556 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_93
timestamp 1666464484
transform 1 0 9660 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_98
timestamp 1666464484
transform 1 0 10120 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_110
timestamp 1666464484
transform 1 0 11224 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_122
timestamp 1666464484
transform 1 0 12328 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_134
timestamp 1666464484
transform 1 0 13432 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_146
timestamp 1666464484
transform 1 0 14536 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_158
timestamp 1666464484
transform 1 0 15640 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_163
timestamp 1666464484
transform 1 0 16100 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_175
timestamp 1666464484
transform 1 0 17204 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_187
timestamp 1666464484
transform 1 0 18308 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_199
timestamp 1666464484
transform 1 0 19412 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_211
timestamp 1666464484
transform 1 0 20516 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_223
timestamp 1666464484
transform 1 0 21620 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_228
timestamp 1666464484
transform 1 0 22080 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_240
timestamp 1666464484
transform 1 0 23184 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_252
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_264
timestamp 1666464484
transform 1 0 25392 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_276
timestamp 1666464484
transform 1 0 26496 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_288
timestamp 1666464484
transform 1 0 27600 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_293
timestamp 1666464484
transform 1 0 28060 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_305
timestamp 1666464484
transform 1 0 29164 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_317
timestamp 1666464484
transform 1 0 30268 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_329
timestamp 1666464484
transform 1 0 31372 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_341
timestamp 1666464484
transform 1 0 32476 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_353
timestamp 1666464484
transform 1 0 33580 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_358
timestamp 1666464484
transform 1 0 34040 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_370
timestamp 1666464484
transform 1 0 35144 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_382
timestamp 1666464484
transform 1 0 36248 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_394
timestamp 1666464484
transform 1 0 37352 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_406
timestamp 1666464484
transform 1 0 38456 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_418
timestamp 1666464484
transform 1 0 39560 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_423
timestamp 1666464484
transform 1 0 40020 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_435
timestamp 1666464484
transform 1 0 41124 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_447
timestamp 1666464484
transform 1 0 42228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_459
timestamp 1666464484
transform 1 0 43332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_471
timestamp 1666464484
transform 1 0 44436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_483
timestamp 1666464484
transform 1 0 45540 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_488
timestamp 1666464484
transform 1 0 46000 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_500
timestamp 1666464484
transform 1 0 47104 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_512
timestamp 1666464484
transform 1 0 48208 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_524
timestamp 1666464484
transform 1 0 49312 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_536
timestamp 1666464484
transform 1 0 50416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_548
timestamp 1666464484
transform 1 0 51520 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_553
timestamp 1666464484
transform 1 0 51980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_565
timestamp 1666464484
transform 1 0 53084 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_577
timestamp 1666464484
transform 1 0 54188 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1666464484
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1666464484
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_613
timestamp 1666464484
transform 1 0 57500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_618
timestamp 1666464484
transform 1 0 57960 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_624
timestamp 1666464484
transform 1 0 58512 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_51
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_63
timestamp 1666464484
transform 1 0 6900 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_66
timestamp 1666464484
transform 1 0 7176 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_78
timestamp 1666464484
transform 1 0 8280 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_90
timestamp 1666464484
transform 1 0 9384 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_102
timestamp 1666464484
transform 1 0 10488 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_114
timestamp 1666464484
transform 1 0 11592 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_126
timestamp 1666464484
transform 1 0 12696 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_131
timestamp 1666464484
transform 1 0 13156 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_143
timestamp 1666464484
transform 1 0 14260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_155
timestamp 1666464484
transform 1 0 15364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_179
timestamp 1666464484
transform 1 0 17572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_191
timestamp 1666464484
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_196
timestamp 1666464484
transform 1 0 19136 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_208
timestamp 1666464484
transform 1 0 20240 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_220
timestamp 1666464484
transform 1 0 21344 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_232
timestamp 1666464484
transform 1 0 22448 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_244
timestamp 1666464484
transform 1 0 23552 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_256
timestamp 1666464484
transform 1 0 24656 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1666464484
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_273
timestamp 1666464484
transform 1 0 26220 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_285
timestamp 1666464484
transform 1 0 27324 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_297
timestamp 1666464484
transform 1 0 28428 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_309
timestamp 1666464484
transform 1 0 29532 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_321
timestamp 1666464484
transform 1 0 30636 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_326
timestamp 1666464484
transform 1 0 31096 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_338
timestamp 1666464484
transform 1 0 32200 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_350
timestamp 1666464484
transform 1 0 33304 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_362
timestamp 1666464484
transform 1 0 34408 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_374
timestamp 1666464484
transform 1 0 35512 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_386
timestamp 1666464484
transform 1 0 36616 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_391
timestamp 1666464484
transform 1 0 37076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_403
timestamp 1666464484
transform 1 0 38180 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_415
timestamp 1666464484
transform 1 0 39284 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_427
timestamp 1666464484
transform 1 0 40388 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_439
timestamp 1666464484
transform 1 0 41492 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_451
timestamp 1666464484
transform 1 0 42596 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_456
timestamp 1666464484
transform 1 0 43056 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_468
timestamp 1666464484
transform 1 0 44160 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_480
timestamp 1666464484
transform 1 0 45264 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_492
timestamp 1666464484
transform 1 0 46368 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_504
timestamp 1666464484
transform 1 0 47472 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_516
timestamp 1666464484
transform 1 0 48576 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_521
timestamp 1666464484
transform 1 0 49036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_533
timestamp 1666464484
transform 1 0 50140 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_545
timestamp 1666464484
transform 1 0 51244 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_557
timestamp 1666464484
transform 1 0 52348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_569
timestamp 1666464484
transform 1 0 53452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_581
timestamp 1666464484
transform 1 0 54556 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_586
timestamp 1666464484
transform 1 0 55016 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_598
timestamp 1666464484
transform 1 0 56120 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_610
timestamp 1666464484
transform 1 0 57224 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_622
timestamp 1666464484
transform 1 0 58328 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_31
timestamp 1666464484
transform 1 0 3956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_33
timestamp 1666464484
transform 1 0 4140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_45
timestamp 1666464484
transform 1 0 5244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_57
timestamp 1666464484
transform 1 0 6348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_69
timestamp 1666464484
transform 1 0 7452 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_81
timestamp 1666464484
transform 1 0 8556 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1666464484
transform 1 0 9660 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_98
timestamp 1666464484
transform 1 0 10120 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_110
timestamp 1666464484
transform 1 0 11224 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_122
timestamp 1666464484
transform 1 0 12328 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_134
timestamp 1666464484
transform 1 0 13432 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_146
timestamp 1666464484
transform 1 0 14536 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_158
timestamp 1666464484
transform 1 0 15640 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_163
timestamp 1666464484
transform 1 0 16100 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_175
timestamp 1666464484
transform 1 0 17204 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_187
timestamp 1666464484
transform 1 0 18308 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_199
timestamp 1666464484
transform 1 0 19412 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_211
timestamp 1666464484
transform 1 0 20516 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_223
timestamp 1666464484
transform 1 0 21620 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_228
timestamp 1666464484
transform 1 0 22080 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_240
timestamp 1666464484
transform 1 0 23184 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_252
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_264
timestamp 1666464484
transform 1 0 25392 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_276
timestamp 1666464484
transform 1 0 26496 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_288
timestamp 1666464484
transform 1 0 27600 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_293
timestamp 1666464484
transform 1 0 28060 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_305
timestamp 1666464484
transform 1 0 29164 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_317
timestamp 1666464484
transform 1 0 30268 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_329
timestamp 1666464484
transform 1 0 31372 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_341
timestamp 1666464484
transform 1 0 32476 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_353
timestamp 1666464484
transform 1 0 33580 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_358
timestamp 1666464484
transform 1 0 34040 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_370
timestamp 1666464484
transform 1 0 35144 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_382
timestamp 1666464484
transform 1 0 36248 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_394
timestamp 1666464484
transform 1 0 37352 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_406
timestamp 1666464484
transform 1 0 38456 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_418
timestamp 1666464484
transform 1 0 39560 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_423
timestamp 1666464484
transform 1 0 40020 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_435
timestamp 1666464484
transform 1 0 41124 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_447
timestamp 1666464484
transform 1 0 42228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_459
timestamp 1666464484
transform 1 0 43332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_471
timestamp 1666464484
transform 1 0 44436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_483
timestamp 1666464484
transform 1 0 45540 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_488
timestamp 1666464484
transform 1 0 46000 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_500
timestamp 1666464484
transform 1 0 47104 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_512
timestamp 1666464484
transform 1 0 48208 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_524
timestamp 1666464484
transform 1 0 49312 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_536
timestamp 1666464484
transform 1 0 50416 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_548
timestamp 1666464484
transform 1 0 51520 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_553
timestamp 1666464484
transform 1 0 51980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_565
timestamp 1666464484
transform 1 0 53084 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_577
timestamp 1666464484
transform 1 0 54188 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1666464484
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1666464484
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_613
timestamp 1666464484
transform 1 0 57500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_618
timestamp 1666464484
transform 1 0 57960 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_624
timestamp 1666464484
transform 1 0 58512 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666464484
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_51
timestamp 1666464484
transform 1 0 5796 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_63
timestamp 1666464484
transform 1 0 6900 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_66
timestamp 1666464484
transform 1 0 7176 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_78
timestamp 1666464484
transform 1 0 8280 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_90
timestamp 1666464484
transform 1 0 9384 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_102
timestamp 1666464484
transform 1 0 10488 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_114
timestamp 1666464484
transform 1 0 11592 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_126
timestamp 1666464484
transform 1 0 12696 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_131
timestamp 1666464484
transform 1 0 13156 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_143
timestamp 1666464484
transform 1 0 14260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_155
timestamp 1666464484
transform 1 0 15364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_179
timestamp 1666464484
transform 1 0 17572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1666464484
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_196
timestamp 1666464484
transform 1 0 19136 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_208
timestamp 1666464484
transform 1 0 20240 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_220
timestamp 1666464484
transform 1 0 21344 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_232
timestamp 1666464484
transform 1 0 22448 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_244
timestamp 1666464484
transform 1 0 23552 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_256
timestamp 1666464484
transform 1 0 24656 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1666464484
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_273
timestamp 1666464484
transform 1 0 26220 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_285
timestamp 1666464484
transform 1 0 27324 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_297
timestamp 1666464484
transform 1 0 28428 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_309
timestamp 1666464484
transform 1 0 29532 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_321
timestamp 1666464484
transform 1 0 30636 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_326
timestamp 1666464484
transform 1 0 31096 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_338
timestamp 1666464484
transform 1 0 32200 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_350
timestamp 1666464484
transform 1 0 33304 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_362
timestamp 1666464484
transform 1 0 34408 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_374
timestamp 1666464484
transform 1 0 35512 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_386
timestamp 1666464484
transform 1 0 36616 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_391
timestamp 1666464484
transform 1 0 37076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_403
timestamp 1666464484
transform 1 0 38180 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_415
timestamp 1666464484
transform 1 0 39284 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_427
timestamp 1666464484
transform 1 0 40388 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_439
timestamp 1666464484
transform 1 0 41492 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_451
timestamp 1666464484
transform 1 0 42596 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_456
timestamp 1666464484
transform 1 0 43056 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_468
timestamp 1666464484
transform 1 0 44160 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_480
timestamp 1666464484
transform 1 0 45264 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_492
timestamp 1666464484
transform 1 0 46368 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_504
timestamp 1666464484
transform 1 0 47472 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_516
timestamp 1666464484
transform 1 0 48576 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_521
timestamp 1666464484
transform 1 0 49036 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_533
timestamp 1666464484
transform 1 0 50140 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_545
timestamp 1666464484
transform 1 0 51244 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_557
timestamp 1666464484
transform 1 0 52348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_569
timestamp 1666464484
transform 1 0 53452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_581
timestamp 1666464484
transform 1 0 54556 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_586
timestamp 1666464484
transform 1 0 55016 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_598
timestamp 1666464484
transform 1 0 56120 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_610
timestamp 1666464484
transform 1 0 57224 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_622
timestamp 1666464484
transform 1 0 58328 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_31
timestamp 1666464484
transform 1 0 3956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_33
timestamp 1666464484
transform 1 0 4140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_45
timestamp 1666464484
transform 1 0 5244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_57
timestamp 1666464484
transform 1 0 6348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_69
timestamp 1666464484
transform 1 0 7452 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_81
timestamp 1666464484
transform 1 0 8556 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_93
timestamp 1666464484
transform 1 0 9660 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_98
timestamp 1666464484
transform 1 0 10120 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_110
timestamp 1666464484
transform 1 0 11224 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_122
timestamp 1666464484
transform 1 0 12328 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_134
timestamp 1666464484
transform 1 0 13432 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_146
timestamp 1666464484
transform 1 0 14536 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_158
timestamp 1666464484
transform 1 0 15640 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_163
timestamp 1666464484
transform 1 0 16100 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_175
timestamp 1666464484
transform 1 0 17204 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_187
timestamp 1666464484
transform 1 0 18308 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_199
timestamp 1666464484
transform 1 0 19412 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_211
timestamp 1666464484
transform 1 0 20516 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_223
timestamp 1666464484
transform 1 0 21620 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_228
timestamp 1666464484
transform 1 0 22080 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_240
timestamp 1666464484
transform 1 0 23184 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_252
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_264
timestamp 1666464484
transform 1 0 25392 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_276
timestamp 1666464484
transform 1 0 26496 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_288
timestamp 1666464484
transform 1 0 27600 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_293
timestamp 1666464484
transform 1 0 28060 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_305
timestamp 1666464484
transform 1 0 29164 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_317
timestamp 1666464484
transform 1 0 30268 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_329
timestamp 1666464484
transform 1 0 31372 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_341
timestamp 1666464484
transform 1 0 32476 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_353
timestamp 1666464484
transform 1 0 33580 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_358
timestamp 1666464484
transform 1 0 34040 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_370
timestamp 1666464484
transform 1 0 35144 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_382
timestamp 1666464484
transform 1 0 36248 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_394
timestamp 1666464484
transform 1 0 37352 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_406
timestamp 1666464484
transform 1 0 38456 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_418
timestamp 1666464484
transform 1 0 39560 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_423
timestamp 1666464484
transform 1 0 40020 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_435
timestamp 1666464484
transform 1 0 41124 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_447
timestamp 1666464484
transform 1 0 42228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_459
timestamp 1666464484
transform 1 0 43332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_471
timestamp 1666464484
transform 1 0 44436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_483
timestamp 1666464484
transform 1 0 45540 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_488
timestamp 1666464484
transform 1 0 46000 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_500
timestamp 1666464484
transform 1 0 47104 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_512
timestamp 1666464484
transform 1 0 48208 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_524
timestamp 1666464484
transform 1 0 49312 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_536
timestamp 1666464484
transform 1 0 50416 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_548
timestamp 1666464484
transform 1 0 51520 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_553
timestamp 1666464484
transform 1 0 51980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_565
timestamp 1666464484
transform 1 0 53084 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_577
timestamp 1666464484
transform 1 0 54188 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1666464484
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1666464484
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_613
timestamp 1666464484
transform 1 0 57500 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_618
timestamp 1666464484
transform 1 0 57960 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_624
timestamp 1666464484
transform 1 0 58512 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1666464484
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_51
timestamp 1666464484
transform 1 0 5796 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_63
timestamp 1666464484
transform 1 0 6900 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_66
timestamp 1666464484
transform 1 0 7176 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_78
timestamp 1666464484
transform 1 0 8280 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_90
timestamp 1666464484
transform 1 0 9384 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_102
timestamp 1666464484
transform 1 0 10488 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_114
timestamp 1666464484
transform 1 0 11592 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_126
timestamp 1666464484
transform 1 0 12696 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_131
timestamp 1666464484
transform 1 0 13156 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_143
timestamp 1666464484
transform 1 0 14260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_155
timestamp 1666464484
transform 1 0 15364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_179
timestamp 1666464484
transform 1 0 17572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_191
timestamp 1666464484
transform 1 0 18676 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_196
timestamp 1666464484
transform 1 0 19136 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_208
timestamp 1666464484
transform 1 0 20240 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_220
timestamp 1666464484
transform 1 0 21344 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_232
timestamp 1666464484
transform 1 0 22448 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_244
timestamp 1666464484
transform 1 0 23552 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_256
timestamp 1666464484
transform 1 0 24656 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1666464484
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_273
timestamp 1666464484
transform 1 0 26220 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_285
timestamp 1666464484
transform 1 0 27324 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_297
timestamp 1666464484
transform 1 0 28428 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_309
timestamp 1666464484
transform 1 0 29532 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_321
timestamp 1666464484
transform 1 0 30636 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_326
timestamp 1666464484
transform 1 0 31096 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_338
timestamp 1666464484
transform 1 0 32200 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_350
timestamp 1666464484
transform 1 0 33304 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_362
timestamp 1666464484
transform 1 0 34408 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_374
timestamp 1666464484
transform 1 0 35512 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_386
timestamp 1666464484
transform 1 0 36616 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_391
timestamp 1666464484
transform 1 0 37076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_403
timestamp 1666464484
transform 1 0 38180 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_415
timestamp 1666464484
transform 1 0 39284 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_427
timestamp 1666464484
transform 1 0 40388 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_439
timestamp 1666464484
transform 1 0 41492 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_451
timestamp 1666464484
transform 1 0 42596 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_456
timestamp 1666464484
transform 1 0 43056 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_468
timestamp 1666464484
transform 1 0 44160 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_480
timestamp 1666464484
transform 1 0 45264 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_492
timestamp 1666464484
transform 1 0 46368 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_504
timestamp 1666464484
transform 1 0 47472 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_516
timestamp 1666464484
transform 1 0 48576 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_521
timestamp 1666464484
transform 1 0 49036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_533
timestamp 1666464484
transform 1 0 50140 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_545
timestamp 1666464484
transform 1 0 51244 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_557
timestamp 1666464484
transform 1 0 52348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_569
timestamp 1666464484
transform 1 0 53452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_581
timestamp 1666464484
transform 1 0 54556 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_586
timestamp 1666464484
transform 1 0 55016 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_598
timestamp 1666464484
transform 1 0 56120 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_610
timestamp 1666464484
transform 1 0 57224 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_622
timestamp 1666464484
transform 1 0 58328 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_31
timestamp 1666464484
transform 1 0 3956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_33
timestamp 1666464484
transform 1 0 4140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_45
timestamp 1666464484
transform 1 0 5244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_57
timestamp 1666464484
transform 1 0 6348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_69
timestamp 1666464484
transform 1 0 7452 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_81
timestamp 1666464484
transform 1 0 8556 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_93
timestamp 1666464484
transform 1 0 9660 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_98
timestamp 1666464484
transform 1 0 10120 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_110
timestamp 1666464484
transform 1 0 11224 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_122
timestamp 1666464484
transform 1 0 12328 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_134
timestamp 1666464484
transform 1 0 13432 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_146
timestamp 1666464484
transform 1 0 14536 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_158
timestamp 1666464484
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_163
timestamp 1666464484
transform 1 0 16100 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_175
timestamp 1666464484
transform 1 0 17204 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_187
timestamp 1666464484
transform 1 0 18308 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_199
timestamp 1666464484
transform 1 0 19412 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_211
timestamp 1666464484
transform 1 0 20516 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_223
timestamp 1666464484
transform 1 0 21620 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_228
timestamp 1666464484
transform 1 0 22080 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_240
timestamp 1666464484
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_252
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_264
timestamp 1666464484
transform 1 0 25392 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_276
timestamp 1666464484
transform 1 0 26496 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1666464484
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_293
timestamp 1666464484
transform 1 0 28060 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_305
timestamp 1666464484
transform 1 0 29164 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_317
timestamp 1666464484
transform 1 0 30268 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_329
timestamp 1666464484
transform 1 0 31372 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_341
timestamp 1666464484
transform 1 0 32476 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_353
timestamp 1666464484
transform 1 0 33580 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_358
timestamp 1666464484
transform 1 0 34040 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_370
timestamp 1666464484
transform 1 0 35144 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_382
timestamp 1666464484
transform 1 0 36248 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_394
timestamp 1666464484
transform 1 0 37352 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_406
timestamp 1666464484
transform 1 0 38456 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_418
timestamp 1666464484
transform 1 0 39560 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_423
timestamp 1666464484
transform 1 0 40020 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_435
timestamp 1666464484
transform 1 0 41124 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_447
timestamp 1666464484
transform 1 0 42228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_459
timestamp 1666464484
transform 1 0 43332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_471
timestamp 1666464484
transform 1 0 44436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_483
timestamp 1666464484
transform 1 0 45540 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_488
timestamp 1666464484
transform 1 0 46000 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_500
timestamp 1666464484
transform 1 0 47104 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_512
timestamp 1666464484
transform 1 0 48208 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_524
timestamp 1666464484
transform 1 0 49312 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_536
timestamp 1666464484
transform 1 0 50416 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_548
timestamp 1666464484
transform 1 0 51520 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_553
timestamp 1666464484
transform 1 0 51980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_565
timestamp 1666464484
transform 1 0 53084 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_577
timestamp 1666464484
transform 1 0 54188 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1666464484
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1666464484
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_613
timestamp 1666464484
transform 1 0 57500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_618
timestamp 1666464484
transform 1 0 57960 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_624
timestamp 1666464484
transform 1 0 58512 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666464484
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1666464484
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1666464484
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_51
timestamp 1666464484
transform 1 0 5796 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_63
timestamp 1666464484
transform 1 0 6900 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_66
timestamp 1666464484
transform 1 0 7176 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_78
timestamp 1666464484
transform 1 0 8280 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_90
timestamp 1666464484
transform 1 0 9384 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_102
timestamp 1666464484
transform 1 0 10488 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_114
timestamp 1666464484
transform 1 0 11592 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_126
timestamp 1666464484
transform 1 0 12696 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_131
timestamp 1666464484
transform 1 0 13156 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_143
timestamp 1666464484
transform 1 0 14260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_155
timestamp 1666464484
transform 1 0 15364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_179
timestamp 1666464484
transform 1 0 17572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1666464484
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_196
timestamp 1666464484
transform 1 0 19136 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_208
timestamp 1666464484
transform 1 0 20240 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_220
timestamp 1666464484
transform 1 0 21344 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_232
timestamp 1666464484
transform 1 0 22448 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_244
timestamp 1666464484
transform 1 0 23552 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_256
timestamp 1666464484
transform 1 0 24656 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1666464484
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_273
timestamp 1666464484
transform 1 0 26220 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_285
timestamp 1666464484
transform 1 0 27324 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_297
timestamp 1666464484
transform 1 0 28428 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_309
timestamp 1666464484
transform 1 0 29532 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_321
timestamp 1666464484
transform 1 0 30636 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_326
timestamp 1666464484
transform 1 0 31096 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_338
timestamp 1666464484
transform 1 0 32200 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_350
timestamp 1666464484
transform 1 0 33304 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_362
timestamp 1666464484
transform 1 0 34408 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_374
timestamp 1666464484
transform 1 0 35512 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_386
timestamp 1666464484
transform 1 0 36616 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_391
timestamp 1666464484
transform 1 0 37076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_403
timestamp 1666464484
transform 1 0 38180 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_415
timestamp 1666464484
transform 1 0 39284 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_427
timestamp 1666464484
transform 1 0 40388 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_439
timestamp 1666464484
transform 1 0 41492 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_451
timestamp 1666464484
transform 1 0 42596 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_456
timestamp 1666464484
transform 1 0 43056 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_468
timestamp 1666464484
transform 1 0 44160 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_480
timestamp 1666464484
transform 1 0 45264 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_492
timestamp 1666464484
transform 1 0 46368 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_504
timestamp 1666464484
transform 1 0 47472 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_516
timestamp 1666464484
transform 1 0 48576 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_521
timestamp 1666464484
transform 1 0 49036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_533
timestamp 1666464484
transform 1 0 50140 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_545
timestamp 1666464484
transform 1 0 51244 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_557
timestamp 1666464484
transform 1 0 52348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_569
timestamp 1666464484
transform 1 0 53452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_581
timestamp 1666464484
transform 1 0 54556 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_586
timestamp 1666464484
transform 1 0 55016 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_598
timestamp 1666464484
transform 1 0 56120 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_610
timestamp 1666464484
transform 1 0 57224 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_622
timestamp 1666464484
transform 1 0 58328 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_31
timestamp 1666464484
transform 1 0 3956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_33
timestamp 1666464484
transform 1 0 4140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_45
timestamp 1666464484
transform 1 0 5244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_57
timestamp 1666464484
transform 1 0 6348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_69
timestamp 1666464484
transform 1 0 7452 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_81
timestamp 1666464484
transform 1 0 8556 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_93
timestamp 1666464484
transform 1 0 9660 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_98
timestamp 1666464484
transform 1 0 10120 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_110
timestamp 1666464484
transform 1 0 11224 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_122
timestamp 1666464484
transform 1 0 12328 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_134
timestamp 1666464484
transform 1 0 13432 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_146
timestamp 1666464484
transform 1 0 14536 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_158
timestamp 1666464484
transform 1 0 15640 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_163
timestamp 1666464484
transform 1 0 16100 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_175
timestamp 1666464484
transform 1 0 17204 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_187
timestamp 1666464484
transform 1 0 18308 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_199
timestamp 1666464484
transform 1 0 19412 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_211
timestamp 1666464484
transform 1 0 20516 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_223
timestamp 1666464484
transform 1 0 21620 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_228
timestamp 1666464484
transform 1 0 22080 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_240
timestamp 1666464484
transform 1 0 23184 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_252
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_264
timestamp 1666464484
transform 1 0 25392 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_276
timestamp 1666464484
transform 1 0 26496 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_288
timestamp 1666464484
transform 1 0 27600 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_293
timestamp 1666464484
transform 1 0 28060 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_305
timestamp 1666464484
transform 1 0 29164 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_317
timestamp 1666464484
transform 1 0 30268 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_329
timestamp 1666464484
transform 1 0 31372 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_341
timestamp 1666464484
transform 1 0 32476 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_353
timestamp 1666464484
transform 1 0 33580 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_358
timestamp 1666464484
transform 1 0 34040 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_370
timestamp 1666464484
transform 1 0 35144 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_382
timestamp 1666464484
transform 1 0 36248 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_394
timestamp 1666464484
transform 1 0 37352 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_406
timestamp 1666464484
transform 1 0 38456 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_418
timestamp 1666464484
transform 1 0 39560 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_423
timestamp 1666464484
transform 1 0 40020 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_435
timestamp 1666464484
transform 1 0 41124 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_447
timestamp 1666464484
transform 1 0 42228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_459
timestamp 1666464484
transform 1 0 43332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_471
timestamp 1666464484
transform 1 0 44436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_483
timestamp 1666464484
transform 1 0 45540 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_488
timestamp 1666464484
transform 1 0 46000 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_500
timestamp 1666464484
transform 1 0 47104 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_512
timestamp 1666464484
transform 1 0 48208 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_524
timestamp 1666464484
transform 1 0 49312 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_536
timestamp 1666464484
transform 1 0 50416 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_548
timestamp 1666464484
transform 1 0 51520 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_553
timestamp 1666464484
transform 1 0 51980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_565
timestamp 1666464484
transform 1 0 53084 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_577
timestamp 1666464484
transform 1 0 54188 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1666464484
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1666464484
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_613
timestamp 1666464484
transform 1 0 57500 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_618
timestamp 1666464484
transform 1 0 57960 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_624
timestamp 1666464484
transform 1 0 58512 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666464484
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666464484
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1666464484
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_51
timestamp 1666464484
transform 1 0 5796 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_63
timestamp 1666464484
transform 1 0 6900 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_66
timestamp 1666464484
transform 1 0 7176 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_78
timestamp 1666464484
transform 1 0 8280 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_90
timestamp 1666464484
transform 1 0 9384 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_102
timestamp 1666464484
transform 1 0 10488 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_114
timestamp 1666464484
transform 1 0 11592 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1666464484
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_131
timestamp 1666464484
transform 1 0 13156 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_143
timestamp 1666464484
transform 1 0 14260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_155
timestamp 1666464484
transform 1 0 15364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_179
timestamp 1666464484
transform 1 0 17572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_191
timestamp 1666464484
transform 1 0 18676 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_196
timestamp 1666464484
transform 1 0 19136 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_208
timestamp 1666464484
transform 1 0 20240 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_220
timestamp 1666464484
transform 1 0 21344 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_232
timestamp 1666464484
transform 1 0 22448 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_244
timestamp 1666464484
transform 1 0 23552 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_256
timestamp 1666464484
transform 1 0 24656 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1666464484
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_273
timestamp 1666464484
transform 1 0 26220 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_285
timestamp 1666464484
transform 1 0 27324 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_297
timestamp 1666464484
transform 1 0 28428 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_309
timestamp 1666464484
transform 1 0 29532 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_321
timestamp 1666464484
transform 1 0 30636 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_326
timestamp 1666464484
transform 1 0 31096 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_338
timestamp 1666464484
transform 1 0 32200 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_350
timestamp 1666464484
transform 1 0 33304 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_362
timestamp 1666464484
transform 1 0 34408 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_374
timestamp 1666464484
transform 1 0 35512 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_386
timestamp 1666464484
transform 1 0 36616 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_391
timestamp 1666464484
transform 1 0 37076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_403
timestamp 1666464484
transform 1 0 38180 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_415
timestamp 1666464484
transform 1 0 39284 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_427
timestamp 1666464484
transform 1 0 40388 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_439
timestamp 1666464484
transform 1 0 41492 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_451
timestamp 1666464484
transform 1 0 42596 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_456
timestamp 1666464484
transform 1 0 43056 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_468
timestamp 1666464484
transform 1 0 44160 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_480
timestamp 1666464484
transform 1 0 45264 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_492
timestamp 1666464484
transform 1 0 46368 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_504
timestamp 1666464484
transform 1 0 47472 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_516
timestamp 1666464484
transform 1 0 48576 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_521
timestamp 1666464484
transform 1 0 49036 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_533
timestamp 1666464484
transform 1 0 50140 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_545
timestamp 1666464484
transform 1 0 51244 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_557
timestamp 1666464484
transform 1 0 52348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_569
timestamp 1666464484
transform 1 0 53452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_581
timestamp 1666464484
transform 1 0 54556 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_586
timestamp 1666464484
transform 1 0 55016 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_598
timestamp 1666464484
transform 1 0 56120 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_610
timestamp 1666464484
transform 1 0 57224 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_622
timestamp 1666464484
transform 1 0 58328 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666464484
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1666464484
transform 1 0 3588 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_31
timestamp 1666464484
transform 1 0 3956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_33
timestamp 1666464484
transform 1 0 4140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_45
timestamp 1666464484
transform 1 0 5244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_57
timestamp 1666464484
transform 1 0 6348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_69
timestamp 1666464484
transform 1 0 7452 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_81
timestamp 1666464484
transform 1 0 8556 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_93
timestamp 1666464484
transform 1 0 9660 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_98
timestamp 1666464484
transform 1 0 10120 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_110
timestamp 1666464484
transform 1 0 11224 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_122
timestamp 1666464484
transform 1 0 12328 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_134
timestamp 1666464484
transform 1 0 13432 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_146
timestamp 1666464484
transform 1 0 14536 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_158
timestamp 1666464484
transform 1 0 15640 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_163
timestamp 1666464484
transform 1 0 16100 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_175
timestamp 1666464484
transform 1 0 17204 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_187
timestamp 1666464484
transform 1 0 18308 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_199
timestamp 1666464484
transform 1 0 19412 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_211
timestamp 1666464484
transform 1 0 20516 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_223
timestamp 1666464484
transform 1 0 21620 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_228
timestamp 1666464484
transform 1 0 22080 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_240
timestamp 1666464484
transform 1 0 23184 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_252
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_264
timestamp 1666464484
transform 1 0 25392 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_276
timestamp 1666464484
transform 1 0 26496 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_288
timestamp 1666464484
transform 1 0 27600 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_293
timestamp 1666464484
transform 1 0 28060 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_305
timestamp 1666464484
transform 1 0 29164 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_317
timestamp 1666464484
transform 1 0 30268 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_329
timestamp 1666464484
transform 1 0 31372 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_341
timestamp 1666464484
transform 1 0 32476 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_353
timestamp 1666464484
transform 1 0 33580 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_358
timestamp 1666464484
transform 1 0 34040 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_370
timestamp 1666464484
transform 1 0 35144 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_382
timestamp 1666464484
transform 1 0 36248 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_394
timestamp 1666464484
transform 1 0 37352 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_406
timestamp 1666464484
transform 1 0 38456 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_418
timestamp 1666464484
transform 1 0 39560 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_423
timestamp 1666464484
transform 1 0 40020 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_435
timestamp 1666464484
transform 1 0 41124 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_447
timestamp 1666464484
transform 1 0 42228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_459
timestamp 1666464484
transform 1 0 43332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_471
timestamp 1666464484
transform 1 0 44436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_483
timestamp 1666464484
transform 1 0 45540 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_488
timestamp 1666464484
transform 1 0 46000 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_500
timestamp 1666464484
transform 1 0 47104 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_512
timestamp 1666464484
transform 1 0 48208 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_524
timestamp 1666464484
transform 1 0 49312 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_536
timestamp 1666464484
transform 1 0 50416 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_548
timestamp 1666464484
transform 1 0 51520 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_553
timestamp 1666464484
transform 1 0 51980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_565
timestamp 1666464484
transform 1 0 53084 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_577
timestamp 1666464484
transform 1 0 54188 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1666464484
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1666464484
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_613
timestamp 1666464484
transform 1 0 57500 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_618
timestamp 1666464484
transform 1 0 57960 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_624
timestamp 1666464484
transform 1 0 58512 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_63
timestamp 1666464484
transform 1 0 6900 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_66
timestamp 1666464484
transform 1 0 7176 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_78
timestamp 1666464484
transform 1 0 8280 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_90
timestamp 1666464484
transform 1 0 9384 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_102
timestamp 1666464484
transform 1 0 10488 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_114
timestamp 1666464484
transform 1 0 11592 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_126
timestamp 1666464484
transform 1 0 12696 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_131
timestamp 1666464484
transform 1 0 13156 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_143
timestamp 1666464484
transform 1 0 14260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_155
timestamp 1666464484
transform 1 0 15364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_167
timestamp 1666464484
transform 1 0 16468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_179
timestamp 1666464484
transform 1 0 17572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_191
timestamp 1666464484
transform 1 0 18676 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_196
timestamp 1666464484
transform 1 0 19136 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_208
timestamp 1666464484
transform 1 0 20240 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_220
timestamp 1666464484
transform 1 0 21344 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_232
timestamp 1666464484
transform 1 0 22448 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_244
timestamp 1666464484
transform 1 0 23552 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_256
timestamp 1666464484
transform 1 0 24656 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1666464484
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_273
timestamp 1666464484
transform 1 0 26220 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_285
timestamp 1666464484
transform 1 0 27324 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_297
timestamp 1666464484
transform 1 0 28428 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_309
timestamp 1666464484
transform 1 0 29532 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_321
timestamp 1666464484
transform 1 0 30636 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_326
timestamp 1666464484
transform 1 0 31096 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_338
timestamp 1666464484
transform 1 0 32200 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_350
timestamp 1666464484
transform 1 0 33304 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_362
timestamp 1666464484
transform 1 0 34408 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_374
timestamp 1666464484
transform 1 0 35512 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_386
timestamp 1666464484
transform 1 0 36616 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_391
timestamp 1666464484
transform 1 0 37076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_403
timestamp 1666464484
transform 1 0 38180 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_415
timestamp 1666464484
transform 1 0 39284 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_427
timestamp 1666464484
transform 1 0 40388 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_439
timestamp 1666464484
transform 1 0 41492 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_451
timestamp 1666464484
transform 1 0 42596 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_456
timestamp 1666464484
transform 1 0 43056 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_468
timestamp 1666464484
transform 1 0 44160 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_480
timestamp 1666464484
transform 1 0 45264 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_492
timestamp 1666464484
transform 1 0 46368 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_504
timestamp 1666464484
transform 1 0 47472 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_516
timestamp 1666464484
transform 1 0 48576 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_521
timestamp 1666464484
transform 1 0 49036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_533
timestamp 1666464484
transform 1 0 50140 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_545
timestamp 1666464484
transform 1 0 51244 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_557
timestamp 1666464484
transform 1 0 52348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_569
timestamp 1666464484
transform 1 0 53452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_581
timestamp 1666464484
transform 1 0 54556 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_586
timestamp 1666464484
transform 1 0 55016 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_598
timestamp 1666464484
transform 1 0 56120 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_610
timestamp 1666464484
transform 1 0 57224 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_622
timestamp 1666464484
transform 1 0 58328 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1666464484
transform 1 0 3588 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_31
timestamp 1666464484
transform 1 0 3956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_33
timestamp 1666464484
transform 1 0 4140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_45
timestamp 1666464484
transform 1 0 5244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_57
timestamp 1666464484
transform 1 0 6348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_69
timestamp 1666464484
transform 1 0 7452 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_81
timestamp 1666464484
transform 1 0 8556 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_93
timestamp 1666464484
transform 1 0 9660 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_98
timestamp 1666464484
transform 1 0 10120 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_110
timestamp 1666464484
transform 1 0 11224 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_122
timestamp 1666464484
transform 1 0 12328 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_134
timestamp 1666464484
transform 1 0 13432 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_146
timestamp 1666464484
transform 1 0 14536 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_158
timestamp 1666464484
transform 1 0 15640 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_163
timestamp 1666464484
transform 1 0 16100 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_175
timestamp 1666464484
transform 1 0 17204 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_187
timestamp 1666464484
transform 1 0 18308 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_199
timestamp 1666464484
transform 1 0 19412 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_211
timestamp 1666464484
transform 1 0 20516 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_223
timestamp 1666464484
transform 1 0 21620 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_228
timestamp 1666464484
transform 1 0 22080 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_240
timestamp 1666464484
transform 1 0 23184 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_252
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_264
timestamp 1666464484
transform 1 0 25392 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_276
timestamp 1666464484
transform 1 0 26496 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_288
timestamp 1666464484
transform 1 0 27600 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_293
timestamp 1666464484
transform 1 0 28060 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_305
timestamp 1666464484
transform 1 0 29164 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_317
timestamp 1666464484
transform 1 0 30268 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_329
timestamp 1666464484
transform 1 0 31372 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_341
timestamp 1666464484
transform 1 0 32476 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_353
timestamp 1666464484
transform 1 0 33580 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_358
timestamp 1666464484
transform 1 0 34040 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_370
timestamp 1666464484
transform 1 0 35144 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_382
timestamp 1666464484
transform 1 0 36248 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_394
timestamp 1666464484
transform 1 0 37352 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_406
timestamp 1666464484
transform 1 0 38456 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_418
timestamp 1666464484
transform 1 0 39560 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_423
timestamp 1666464484
transform 1 0 40020 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_435
timestamp 1666464484
transform 1 0 41124 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_447
timestamp 1666464484
transform 1 0 42228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_459
timestamp 1666464484
transform 1 0 43332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_471
timestamp 1666464484
transform 1 0 44436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_483
timestamp 1666464484
transform 1 0 45540 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_488
timestamp 1666464484
transform 1 0 46000 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_500
timestamp 1666464484
transform 1 0 47104 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_512
timestamp 1666464484
transform 1 0 48208 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_524
timestamp 1666464484
transform 1 0 49312 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_536
timestamp 1666464484
transform 1 0 50416 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_548
timestamp 1666464484
transform 1 0 51520 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_553
timestamp 1666464484
transform 1 0 51980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_565
timestamp 1666464484
transform 1 0 53084 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_577
timestamp 1666464484
transform 1 0 54188 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1666464484
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1666464484
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_613
timestamp 1666464484
transform 1 0 57500 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_618
timestamp 1666464484
transform 1 0 57960 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_624
timestamp 1666464484
transform 1 0 58512 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666464484
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666464484
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1666464484
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_51
timestamp 1666464484
transform 1 0 5796 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_63
timestamp 1666464484
transform 1 0 6900 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_66
timestamp 1666464484
transform 1 0 7176 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_78
timestamp 1666464484
transform 1 0 8280 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_90
timestamp 1666464484
transform 1 0 9384 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_102
timestamp 1666464484
transform 1 0 10488 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_114
timestamp 1666464484
transform 1 0 11592 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_126
timestamp 1666464484
transform 1 0 12696 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_131
timestamp 1666464484
transform 1 0 13156 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_143
timestamp 1666464484
transform 1 0 14260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_155
timestamp 1666464484
transform 1 0 15364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_167
timestamp 1666464484
transform 1 0 16468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_179
timestamp 1666464484
transform 1 0 17572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_191
timestamp 1666464484
transform 1 0 18676 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_196
timestamp 1666464484
transform 1 0 19136 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_208
timestamp 1666464484
transform 1 0 20240 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_220
timestamp 1666464484
transform 1 0 21344 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_232
timestamp 1666464484
transform 1 0 22448 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_244
timestamp 1666464484
transform 1 0 23552 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_256
timestamp 1666464484
transform 1 0 24656 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_273
timestamp 1666464484
transform 1 0 26220 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_285
timestamp 1666464484
transform 1 0 27324 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_297
timestamp 1666464484
transform 1 0 28428 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_309
timestamp 1666464484
transform 1 0 29532 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_321
timestamp 1666464484
transform 1 0 30636 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_326
timestamp 1666464484
transform 1 0 31096 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_338
timestamp 1666464484
transform 1 0 32200 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_350
timestamp 1666464484
transform 1 0 33304 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_362
timestamp 1666464484
transform 1 0 34408 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_374
timestamp 1666464484
transform 1 0 35512 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_386
timestamp 1666464484
transform 1 0 36616 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_391
timestamp 1666464484
transform 1 0 37076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_403
timestamp 1666464484
transform 1 0 38180 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_415
timestamp 1666464484
transform 1 0 39284 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_427
timestamp 1666464484
transform 1 0 40388 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_439
timestamp 1666464484
transform 1 0 41492 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_451
timestamp 1666464484
transform 1 0 42596 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_456
timestamp 1666464484
transform 1 0 43056 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_468
timestamp 1666464484
transform 1 0 44160 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_480
timestamp 1666464484
transform 1 0 45264 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_492
timestamp 1666464484
transform 1 0 46368 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_504
timestamp 1666464484
transform 1 0 47472 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_516
timestamp 1666464484
transform 1 0 48576 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_521
timestamp 1666464484
transform 1 0 49036 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_533
timestamp 1666464484
transform 1 0 50140 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_545
timestamp 1666464484
transform 1 0 51244 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_557
timestamp 1666464484
transform 1 0 52348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_569
timestamp 1666464484
transform 1 0 53452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_581
timestamp 1666464484
transform 1 0 54556 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_586
timestamp 1666464484
transform 1 0 55016 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_598
timestamp 1666464484
transform 1 0 56120 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_610
timestamp 1666464484
transform 1 0 57224 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_622
timestamp 1666464484
transform 1 0 58328 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_31
timestamp 1666464484
transform 1 0 3956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_33
timestamp 1666464484
transform 1 0 4140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_45
timestamp 1666464484
transform 1 0 5244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_57
timestamp 1666464484
transform 1 0 6348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_69
timestamp 1666464484
transform 1 0 7452 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_81
timestamp 1666464484
transform 1 0 8556 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_93
timestamp 1666464484
transform 1 0 9660 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_98
timestamp 1666464484
transform 1 0 10120 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_110
timestamp 1666464484
transform 1 0 11224 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_122
timestamp 1666464484
transform 1 0 12328 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_134
timestamp 1666464484
transform 1 0 13432 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_146
timestamp 1666464484
transform 1 0 14536 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_158
timestamp 1666464484
transform 1 0 15640 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_163
timestamp 1666464484
transform 1 0 16100 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_175
timestamp 1666464484
transform 1 0 17204 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_187
timestamp 1666464484
transform 1 0 18308 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_199
timestamp 1666464484
transform 1 0 19412 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_211
timestamp 1666464484
transform 1 0 20516 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_223
timestamp 1666464484
transform 1 0 21620 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_228
timestamp 1666464484
transform 1 0 22080 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_240
timestamp 1666464484
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_252
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_264
timestamp 1666464484
transform 1 0 25392 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_276
timestamp 1666464484
transform 1 0 26496 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_288
timestamp 1666464484
transform 1 0 27600 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_293
timestamp 1666464484
transform 1 0 28060 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_305
timestamp 1666464484
transform 1 0 29164 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_317
timestamp 1666464484
transform 1 0 30268 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_329
timestamp 1666464484
transform 1 0 31372 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_341
timestamp 1666464484
transform 1 0 32476 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_353
timestamp 1666464484
transform 1 0 33580 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_358
timestamp 1666464484
transform 1 0 34040 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_370
timestamp 1666464484
transform 1 0 35144 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_382
timestamp 1666464484
transform 1 0 36248 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_394
timestamp 1666464484
transform 1 0 37352 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_406
timestamp 1666464484
transform 1 0 38456 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_418
timestamp 1666464484
transform 1 0 39560 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_423
timestamp 1666464484
transform 1 0 40020 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_435
timestamp 1666464484
transform 1 0 41124 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_447
timestamp 1666464484
transform 1 0 42228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_459
timestamp 1666464484
transform 1 0 43332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_471
timestamp 1666464484
transform 1 0 44436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_483
timestamp 1666464484
transform 1 0 45540 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_488
timestamp 1666464484
transform 1 0 46000 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_500
timestamp 1666464484
transform 1 0 47104 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_512
timestamp 1666464484
transform 1 0 48208 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_524
timestamp 1666464484
transform 1 0 49312 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_536
timestamp 1666464484
transform 1 0 50416 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_548
timestamp 1666464484
transform 1 0 51520 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_553
timestamp 1666464484
transform 1 0 51980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_565
timestamp 1666464484
transform 1 0 53084 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_577
timestamp 1666464484
transform 1 0 54188 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1666464484
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1666464484
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_613
timestamp 1666464484
transform 1 0 57500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_618
timestamp 1666464484
transform 1 0 57960 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_624
timestamp 1666464484
transform 1 0 58512 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_63
timestamp 1666464484
transform 1 0 6900 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_66
timestamp 1666464484
transform 1 0 7176 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_78
timestamp 1666464484
transform 1 0 8280 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_90
timestamp 1666464484
transform 1 0 9384 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_102
timestamp 1666464484
transform 1 0 10488 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_114
timestamp 1666464484
transform 1 0 11592 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_126
timestamp 1666464484
transform 1 0 12696 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_131
timestamp 1666464484
transform 1 0 13156 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_143
timestamp 1666464484
transform 1 0 14260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_155
timestamp 1666464484
transform 1 0 15364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_179
timestamp 1666464484
transform 1 0 17572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_191
timestamp 1666464484
transform 1 0 18676 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_196
timestamp 1666464484
transform 1 0 19136 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_208
timestamp 1666464484
transform 1 0 20240 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_220
timestamp 1666464484
transform 1 0 21344 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_232
timestamp 1666464484
transform 1 0 22448 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_244
timestamp 1666464484
transform 1 0 23552 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_256
timestamp 1666464484
transform 1 0 24656 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1666464484
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_273
timestamp 1666464484
transform 1 0 26220 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_285
timestamp 1666464484
transform 1 0 27324 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_297
timestamp 1666464484
transform 1 0 28428 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_309
timestamp 1666464484
transform 1 0 29532 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_321
timestamp 1666464484
transform 1 0 30636 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_326
timestamp 1666464484
transform 1 0 31096 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_338
timestamp 1666464484
transform 1 0 32200 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_350
timestamp 1666464484
transform 1 0 33304 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_362
timestamp 1666464484
transform 1 0 34408 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_374
timestamp 1666464484
transform 1 0 35512 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_386
timestamp 1666464484
transform 1 0 36616 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_391
timestamp 1666464484
transform 1 0 37076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_403
timestamp 1666464484
transform 1 0 38180 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_415
timestamp 1666464484
transform 1 0 39284 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_427
timestamp 1666464484
transform 1 0 40388 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_439
timestamp 1666464484
transform 1 0 41492 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_451
timestamp 1666464484
transform 1 0 42596 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_456
timestamp 1666464484
transform 1 0 43056 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_468
timestamp 1666464484
transform 1 0 44160 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_480
timestamp 1666464484
transform 1 0 45264 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_492
timestamp 1666464484
transform 1 0 46368 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_504
timestamp 1666464484
transform 1 0 47472 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_516
timestamp 1666464484
transform 1 0 48576 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_521
timestamp 1666464484
transform 1 0 49036 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_533
timestamp 1666464484
transform 1 0 50140 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_545
timestamp 1666464484
transform 1 0 51244 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_557
timestamp 1666464484
transform 1 0 52348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_569
timestamp 1666464484
transform 1 0 53452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_581
timestamp 1666464484
transform 1 0 54556 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_586
timestamp 1666464484
transform 1 0 55016 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_598
timestamp 1666464484
transform 1 0 56120 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_610
timestamp 1666464484
transform 1 0 57224 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_622
timestamp 1666464484
transform 1 0 58328 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_31
timestamp 1666464484
transform 1 0 3956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_33
timestamp 1666464484
transform 1 0 4140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_45
timestamp 1666464484
transform 1 0 5244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_57
timestamp 1666464484
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_69
timestamp 1666464484
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_81
timestamp 1666464484
transform 1 0 8556 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_93
timestamp 1666464484
transform 1 0 9660 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_98
timestamp 1666464484
transform 1 0 10120 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_110
timestamp 1666464484
transform 1 0 11224 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_122
timestamp 1666464484
transform 1 0 12328 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_134
timestamp 1666464484
transform 1 0 13432 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_146
timestamp 1666464484
transform 1 0 14536 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_158
timestamp 1666464484
transform 1 0 15640 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_163
timestamp 1666464484
transform 1 0 16100 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_175
timestamp 1666464484
transform 1 0 17204 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_187
timestamp 1666464484
transform 1 0 18308 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_199
timestamp 1666464484
transform 1 0 19412 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_211
timestamp 1666464484
transform 1 0 20516 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_223
timestamp 1666464484
transform 1 0 21620 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_228
timestamp 1666464484
transform 1 0 22080 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_240
timestamp 1666464484
transform 1 0 23184 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_252
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_264
timestamp 1666464484
transform 1 0 25392 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_276
timestamp 1666464484
transform 1 0 26496 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_288
timestamp 1666464484
transform 1 0 27600 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_293
timestamp 1666464484
transform 1 0 28060 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_305
timestamp 1666464484
transform 1 0 29164 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_317
timestamp 1666464484
transform 1 0 30268 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_329
timestamp 1666464484
transform 1 0 31372 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_341
timestamp 1666464484
transform 1 0 32476 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_353
timestamp 1666464484
transform 1 0 33580 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_358
timestamp 1666464484
transform 1 0 34040 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_370
timestamp 1666464484
transform 1 0 35144 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_382
timestamp 1666464484
transform 1 0 36248 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_394
timestamp 1666464484
transform 1 0 37352 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_406
timestamp 1666464484
transform 1 0 38456 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_418
timestamp 1666464484
transform 1 0 39560 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_423
timestamp 1666464484
transform 1 0 40020 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_435
timestamp 1666464484
transform 1 0 41124 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_447
timestamp 1666464484
transform 1 0 42228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_459
timestamp 1666464484
transform 1 0 43332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_471
timestamp 1666464484
transform 1 0 44436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_483
timestamp 1666464484
transform 1 0 45540 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_488
timestamp 1666464484
transform 1 0 46000 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_500
timestamp 1666464484
transform 1 0 47104 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_512
timestamp 1666464484
transform 1 0 48208 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_524
timestamp 1666464484
transform 1 0 49312 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_536
timestamp 1666464484
transform 1 0 50416 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_548
timestamp 1666464484
transform 1 0 51520 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_553
timestamp 1666464484
transform 1 0 51980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_565
timestamp 1666464484
transform 1 0 53084 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_577
timestamp 1666464484
transform 1 0 54188 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1666464484
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1666464484
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_613
timestamp 1666464484
transform 1 0 57500 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_618
timestamp 1666464484
transform 1 0 57960 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_624
timestamp 1666464484
transform 1 0 58512 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666464484
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_51
timestamp 1666464484
transform 1 0 5796 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_63
timestamp 1666464484
transform 1 0 6900 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_66
timestamp 1666464484
transform 1 0 7176 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_78
timestamp 1666464484
transform 1 0 8280 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_90
timestamp 1666464484
transform 1 0 9384 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_102
timestamp 1666464484
transform 1 0 10488 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_114
timestamp 1666464484
transform 1 0 11592 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_126
timestamp 1666464484
transform 1 0 12696 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_131
timestamp 1666464484
transform 1 0 13156 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_143
timestamp 1666464484
transform 1 0 14260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_155
timestamp 1666464484
transform 1 0 15364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_167
timestamp 1666464484
transform 1 0 16468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_179
timestamp 1666464484
transform 1 0 17572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_191
timestamp 1666464484
transform 1 0 18676 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_196
timestamp 1666464484
transform 1 0 19136 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_208
timestamp 1666464484
transform 1 0 20240 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_220
timestamp 1666464484
transform 1 0 21344 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_232
timestamp 1666464484
transform 1 0 22448 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_244
timestamp 1666464484
transform 1 0 23552 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_256
timestamp 1666464484
transform 1 0 24656 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1666464484
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_273
timestamp 1666464484
transform 1 0 26220 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_285
timestamp 1666464484
transform 1 0 27324 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_297
timestamp 1666464484
transform 1 0 28428 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_309
timestamp 1666464484
transform 1 0 29532 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_321
timestamp 1666464484
transform 1 0 30636 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_326
timestamp 1666464484
transform 1 0 31096 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_338
timestamp 1666464484
transform 1 0 32200 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_350
timestamp 1666464484
transform 1 0 33304 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_362
timestamp 1666464484
transform 1 0 34408 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_374
timestamp 1666464484
transform 1 0 35512 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_386
timestamp 1666464484
transform 1 0 36616 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_391
timestamp 1666464484
transform 1 0 37076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_403
timestamp 1666464484
transform 1 0 38180 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_415
timestamp 1666464484
transform 1 0 39284 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_427
timestamp 1666464484
transform 1 0 40388 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_439
timestamp 1666464484
transform 1 0 41492 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_451
timestamp 1666464484
transform 1 0 42596 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_456
timestamp 1666464484
transform 1 0 43056 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_468
timestamp 1666464484
transform 1 0 44160 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_480
timestamp 1666464484
transform 1 0 45264 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_492
timestamp 1666464484
transform 1 0 46368 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_504
timestamp 1666464484
transform 1 0 47472 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_516
timestamp 1666464484
transform 1 0 48576 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_521
timestamp 1666464484
transform 1 0 49036 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_533
timestamp 1666464484
transform 1 0 50140 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_545
timestamp 1666464484
transform 1 0 51244 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_557
timestamp 1666464484
transform 1 0 52348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_569
timestamp 1666464484
transform 1 0 53452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_581
timestamp 1666464484
transform 1 0 54556 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_586
timestamp 1666464484
transform 1 0 55016 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_598
timestamp 1666464484
transform 1 0 56120 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_610
timestamp 1666464484
transform 1 0 57224 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_622
timestamp 1666464484
transform 1 0 58328 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1666464484
transform 1 0 3588 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_31
timestamp 1666464484
transform 1 0 3956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_33
timestamp 1666464484
transform 1 0 4140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_45
timestamp 1666464484
transform 1 0 5244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_57
timestamp 1666464484
transform 1 0 6348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_69
timestamp 1666464484
transform 1 0 7452 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_81
timestamp 1666464484
transform 1 0 8556 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_93
timestamp 1666464484
transform 1 0 9660 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_98
timestamp 1666464484
transform 1 0 10120 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_110
timestamp 1666464484
transform 1 0 11224 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_122
timestamp 1666464484
transform 1 0 12328 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_134
timestamp 1666464484
transform 1 0 13432 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_146
timestamp 1666464484
transform 1 0 14536 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_158
timestamp 1666464484
transform 1 0 15640 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_163
timestamp 1666464484
transform 1 0 16100 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_175
timestamp 1666464484
transform 1 0 17204 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_187
timestamp 1666464484
transform 1 0 18308 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_199
timestamp 1666464484
transform 1 0 19412 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_211
timestamp 1666464484
transform 1 0 20516 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_223
timestamp 1666464484
transform 1 0 21620 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_228
timestamp 1666464484
transform 1 0 22080 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_240
timestamp 1666464484
transform 1 0 23184 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_252
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_264
timestamp 1666464484
transform 1 0 25392 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_276
timestamp 1666464484
transform 1 0 26496 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_288
timestamp 1666464484
transform 1 0 27600 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_293
timestamp 1666464484
transform 1 0 28060 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_305
timestamp 1666464484
transform 1 0 29164 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_317
timestamp 1666464484
transform 1 0 30268 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_329
timestamp 1666464484
transform 1 0 31372 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_341
timestamp 1666464484
transform 1 0 32476 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_353
timestamp 1666464484
transform 1 0 33580 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_358
timestamp 1666464484
transform 1 0 34040 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_370
timestamp 1666464484
transform 1 0 35144 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_382
timestamp 1666464484
transform 1 0 36248 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_394
timestamp 1666464484
transform 1 0 37352 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_406
timestamp 1666464484
transform 1 0 38456 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_418
timestamp 1666464484
transform 1 0 39560 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_423
timestamp 1666464484
transform 1 0 40020 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_435
timestamp 1666464484
transform 1 0 41124 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_447
timestamp 1666464484
transform 1 0 42228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_459
timestamp 1666464484
transform 1 0 43332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_471
timestamp 1666464484
transform 1 0 44436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_483
timestamp 1666464484
transform 1 0 45540 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_488
timestamp 1666464484
transform 1 0 46000 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_500
timestamp 1666464484
transform 1 0 47104 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_512
timestamp 1666464484
transform 1 0 48208 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_524
timestamp 1666464484
transform 1 0 49312 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_536
timestamp 1666464484
transform 1 0 50416 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_548
timestamp 1666464484
transform 1 0 51520 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_553
timestamp 1666464484
transform 1 0 51980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_565
timestamp 1666464484
transform 1 0 53084 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_577
timestamp 1666464484
transform 1 0 54188 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1666464484
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1666464484
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_613
timestamp 1666464484
transform 1 0 57500 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_618
timestamp 1666464484
transform 1 0 57960 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_624
timestamp 1666464484
transform 1 0 58512 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_63
timestamp 1666464484
transform 1 0 6900 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_66
timestamp 1666464484
transform 1 0 7176 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_78
timestamp 1666464484
transform 1 0 8280 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_90
timestamp 1666464484
transform 1 0 9384 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_102
timestamp 1666464484
transform 1 0 10488 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_114
timestamp 1666464484
transform 1 0 11592 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_126
timestamp 1666464484
transform 1 0 12696 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_131
timestamp 1666464484
transform 1 0 13156 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_143
timestamp 1666464484
transform 1 0 14260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_155
timestamp 1666464484
transform 1 0 15364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_167
timestamp 1666464484
transform 1 0 16468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_179
timestamp 1666464484
transform 1 0 17572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_191
timestamp 1666464484
transform 1 0 18676 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_196
timestamp 1666464484
transform 1 0 19136 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_208
timestamp 1666464484
transform 1 0 20240 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_220
timestamp 1666464484
transform 1 0 21344 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_232
timestamp 1666464484
transform 1 0 22448 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_244
timestamp 1666464484
transform 1 0 23552 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_256
timestamp 1666464484
transform 1 0 24656 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1666464484
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_273
timestamp 1666464484
transform 1 0 26220 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_285
timestamp 1666464484
transform 1 0 27324 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_297
timestamp 1666464484
transform 1 0 28428 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_309
timestamp 1666464484
transform 1 0 29532 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_321
timestamp 1666464484
transform 1 0 30636 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_326
timestamp 1666464484
transform 1 0 31096 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_338
timestamp 1666464484
transform 1 0 32200 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_350
timestamp 1666464484
transform 1 0 33304 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_362
timestamp 1666464484
transform 1 0 34408 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_374
timestamp 1666464484
transform 1 0 35512 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_386
timestamp 1666464484
transform 1 0 36616 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_391
timestamp 1666464484
transform 1 0 37076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_403
timestamp 1666464484
transform 1 0 38180 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_415
timestamp 1666464484
transform 1 0 39284 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_427
timestamp 1666464484
transform 1 0 40388 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_439
timestamp 1666464484
transform 1 0 41492 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_451
timestamp 1666464484
transform 1 0 42596 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_456
timestamp 1666464484
transform 1 0 43056 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_468
timestamp 1666464484
transform 1 0 44160 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_480
timestamp 1666464484
transform 1 0 45264 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_492
timestamp 1666464484
transform 1 0 46368 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_504
timestamp 1666464484
transform 1 0 47472 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_516
timestamp 1666464484
transform 1 0 48576 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_521
timestamp 1666464484
transform 1 0 49036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_533
timestamp 1666464484
transform 1 0 50140 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_545
timestamp 1666464484
transform 1 0 51244 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_557
timestamp 1666464484
transform 1 0 52348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_569
timestamp 1666464484
transform 1 0 53452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_581
timestamp 1666464484
transform 1 0 54556 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_586
timestamp 1666464484
transform 1 0 55016 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_598
timestamp 1666464484
transform 1 0 56120 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_610
timestamp 1666464484
transform 1 0 57224 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_622
timestamp 1666464484
transform 1 0 58328 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_31
timestamp 1666464484
transform 1 0 3956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_33
timestamp 1666464484
transform 1 0 4140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_45
timestamp 1666464484
transform 1 0 5244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_57
timestamp 1666464484
transform 1 0 6348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_69
timestamp 1666464484
transform 1 0 7452 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_81
timestamp 1666464484
transform 1 0 8556 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_93
timestamp 1666464484
transform 1 0 9660 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_98
timestamp 1666464484
transform 1 0 10120 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_110
timestamp 1666464484
transform 1 0 11224 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_122
timestamp 1666464484
transform 1 0 12328 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_134
timestamp 1666464484
transform 1 0 13432 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_146
timestamp 1666464484
transform 1 0 14536 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_158
timestamp 1666464484
transform 1 0 15640 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_163
timestamp 1666464484
transform 1 0 16100 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_175
timestamp 1666464484
transform 1 0 17204 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_187
timestamp 1666464484
transform 1 0 18308 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_199
timestamp 1666464484
transform 1 0 19412 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_211
timestamp 1666464484
transform 1 0 20516 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_223
timestamp 1666464484
transform 1 0 21620 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_228
timestamp 1666464484
transform 1 0 22080 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_240
timestamp 1666464484
transform 1 0 23184 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_252
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_264
timestamp 1666464484
transform 1 0 25392 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_276
timestamp 1666464484
transform 1 0 26496 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_288
timestamp 1666464484
transform 1 0 27600 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_293
timestamp 1666464484
transform 1 0 28060 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_305
timestamp 1666464484
transform 1 0 29164 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_317
timestamp 1666464484
transform 1 0 30268 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_329
timestamp 1666464484
transform 1 0 31372 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_341
timestamp 1666464484
transform 1 0 32476 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_353
timestamp 1666464484
transform 1 0 33580 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_358
timestamp 1666464484
transform 1 0 34040 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_370
timestamp 1666464484
transform 1 0 35144 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_382
timestamp 1666464484
transform 1 0 36248 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_394
timestamp 1666464484
transform 1 0 37352 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_406
timestamp 1666464484
transform 1 0 38456 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_418
timestamp 1666464484
transform 1 0 39560 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_423
timestamp 1666464484
transform 1 0 40020 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_435
timestamp 1666464484
transform 1 0 41124 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_447
timestamp 1666464484
transform 1 0 42228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_459
timestamp 1666464484
transform 1 0 43332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_471
timestamp 1666464484
transform 1 0 44436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_483
timestamp 1666464484
transform 1 0 45540 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_488
timestamp 1666464484
transform 1 0 46000 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_500
timestamp 1666464484
transform 1 0 47104 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_512
timestamp 1666464484
transform 1 0 48208 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_524
timestamp 1666464484
transform 1 0 49312 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_536
timestamp 1666464484
transform 1 0 50416 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_548
timestamp 1666464484
transform 1 0 51520 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_553
timestamp 1666464484
transform 1 0 51980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_565
timestamp 1666464484
transform 1 0 53084 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_577
timestamp 1666464484
transform 1 0 54188 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1666464484
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1666464484
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_613
timestamp 1666464484
transform 1 0 57500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_618
timestamp 1666464484
transform 1 0 57960 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_624
timestamp 1666464484
transform 1 0 58512 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_63
timestamp 1666464484
transform 1 0 6900 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_66
timestamp 1666464484
transform 1 0 7176 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_78
timestamp 1666464484
transform 1 0 8280 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_90
timestamp 1666464484
transform 1 0 9384 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_102
timestamp 1666464484
transform 1 0 10488 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_114
timestamp 1666464484
transform 1 0 11592 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_126
timestamp 1666464484
transform 1 0 12696 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_131
timestamp 1666464484
transform 1 0 13156 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_143
timestamp 1666464484
transform 1 0 14260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_155
timestamp 1666464484
transform 1 0 15364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_167
timestamp 1666464484
transform 1 0 16468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_179
timestamp 1666464484
transform 1 0 17572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_191
timestamp 1666464484
transform 1 0 18676 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_196
timestamp 1666464484
transform 1 0 19136 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_208
timestamp 1666464484
transform 1 0 20240 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_220
timestamp 1666464484
transform 1 0 21344 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_232
timestamp 1666464484
transform 1 0 22448 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_244
timestamp 1666464484
transform 1 0 23552 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_256
timestamp 1666464484
transform 1 0 24656 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1666464484
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_273
timestamp 1666464484
transform 1 0 26220 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_285
timestamp 1666464484
transform 1 0 27324 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_297
timestamp 1666464484
transform 1 0 28428 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_309
timestamp 1666464484
transform 1 0 29532 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_321
timestamp 1666464484
transform 1 0 30636 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_326
timestamp 1666464484
transform 1 0 31096 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_338
timestamp 1666464484
transform 1 0 32200 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_350
timestamp 1666464484
transform 1 0 33304 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_362
timestamp 1666464484
transform 1 0 34408 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_374
timestamp 1666464484
transform 1 0 35512 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_386
timestamp 1666464484
transform 1 0 36616 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_391
timestamp 1666464484
transform 1 0 37076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_403
timestamp 1666464484
transform 1 0 38180 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_415
timestamp 1666464484
transform 1 0 39284 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_427
timestamp 1666464484
transform 1 0 40388 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_439
timestamp 1666464484
transform 1 0 41492 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_451
timestamp 1666464484
transform 1 0 42596 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_456
timestamp 1666464484
transform 1 0 43056 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_468
timestamp 1666464484
transform 1 0 44160 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_480
timestamp 1666464484
transform 1 0 45264 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_492
timestamp 1666464484
transform 1 0 46368 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_504
timestamp 1666464484
transform 1 0 47472 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_516
timestamp 1666464484
transform 1 0 48576 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_521
timestamp 1666464484
transform 1 0 49036 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_533
timestamp 1666464484
transform 1 0 50140 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_545
timestamp 1666464484
transform 1 0 51244 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_557
timestamp 1666464484
transform 1 0 52348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_569
timestamp 1666464484
transform 1 0 53452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_581
timestamp 1666464484
transform 1 0 54556 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_586
timestamp 1666464484
transform 1 0 55016 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_598
timestamp 1666464484
transform 1 0 56120 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_610
timestamp 1666464484
transform 1 0 57224 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_622
timestamp 1666464484
transform 1 0 58328 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_31
timestamp 1666464484
transform 1 0 3956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_33
timestamp 1666464484
transform 1 0 4140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_45
timestamp 1666464484
transform 1 0 5244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_57
timestamp 1666464484
transform 1 0 6348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_69
timestamp 1666464484
transform 1 0 7452 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_81
timestamp 1666464484
transform 1 0 8556 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_93
timestamp 1666464484
transform 1 0 9660 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_98
timestamp 1666464484
transform 1 0 10120 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_110
timestamp 1666464484
transform 1 0 11224 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_122
timestamp 1666464484
transform 1 0 12328 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_134
timestamp 1666464484
transform 1 0 13432 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_146
timestamp 1666464484
transform 1 0 14536 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_158
timestamp 1666464484
transform 1 0 15640 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_163
timestamp 1666464484
transform 1 0 16100 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_175
timestamp 1666464484
transform 1 0 17204 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_187
timestamp 1666464484
transform 1 0 18308 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_199
timestamp 1666464484
transform 1 0 19412 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_211
timestamp 1666464484
transform 1 0 20516 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_223
timestamp 1666464484
transform 1 0 21620 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_228
timestamp 1666464484
transform 1 0 22080 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_240
timestamp 1666464484
transform 1 0 23184 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_252
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_264
timestamp 1666464484
transform 1 0 25392 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_276
timestamp 1666464484
transform 1 0 26496 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_288
timestamp 1666464484
transform 1 0 27600 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_293
timestamp 1666464484
transform 1 0 28060 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_305
timestamp 1666464484
transform 1 0 29164 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_317
timestamp 1666464484
transform 1 0 30268 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_329
timestamp 1666464484
transform 1 0 31372 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_341
timestamp 1666464484
transform 1 0 32476 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_353
timestamp 1666464484
transform 1 0 33580 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_358
timestamp 1666464484
transform 1 0 34040 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_370
timestamp 1666464484
transform 1 0 35144 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_382
timestamp 1666464484
transform 1 0 36248 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_394
timestamp 1666464484
transform 1 0 37352 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_406
timestamp 1666464484
transform 1 0 38456 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_418
timestamp 1666464484
transform 1 0 39560 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_423
timestamp 1666464484
transform 1 0 40020 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_435
timestamp 1666464484
transform 1 0 41124 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_447
timestamp 1666464484
transform 1 0 42228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_459
timestamp 1666464484
transform 1 0 43332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_471
timestamp 1666464484
transform 1 0 44436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_483
timestamp 1666464484
transform 1 0 45540 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_488
timestamp 1666464484
transform 1 0 46000 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_500
timestamp 1666464484
transform 1 0 47104 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_512
timestamp 1666464484
transform 1 0 48208 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_524
timestamp 1666464484
transform 1 0 49312 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_536
timestamp 1666464484
transform 1 0 50416 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_548
timestamp 1666464484
transform 1 0 51520 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_553
timestamp 1666464484
transform 1 0 51980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_565
timestamp 1666464484
transform 1 0 53084 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_577
timestamp 1666464484
transform 1 0 54188 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1666464484
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1666464484
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_613
timestamp 1666464484
transform 1 0 57500 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_618
timestamp 1666464484
transform 1 0 57960 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_624
timestamp 1666464484
transform 1 0 58512 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666464484
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666464484
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1666464484
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_51
timestamp 1666464484
transform 1 0 5796 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_63
timestamp 1666464484
transform 1 0 6900 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_66
timestamp 1666464484
transform 1 0 7176 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_78
timestamp 1666464484
transform 1 0 8280 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_90
timestamp 1666464484
transform 1 0 9384 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_102
timestamp 1666464484
transform 1 0 10488 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_114
timestamp 1666464484
transform 1 0 11592 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_126
timestamp 1666464484
transform 1 0 12696 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_131
timestamp 1666464484
transform 1 0 13156 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_143
timestamp 1666464484
transform 1 0 14260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_155
timestamp 1666464484
transform 1 0 15364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_167
timestamp 1666464484
transform 1 0 16468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_179
timestamp 1666464484
transform 1 0 17572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_191
timestamp 1666464484
transform 1 0 18676 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_196
timestamp 1666464484
transform 1 0 19136 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_208
timestamp 1666464484
transform 1 0 20240 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_220
timestamp 1666464484
transform 1 0 21344 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_232
timestamp 1666464484
transform 1 0 22448 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_244
timestamp 1666464484
transform 1 0 23552 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1666464484
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1666464484
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_273
timestamp 1666464484
transform 1 0 26220 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_285
timestamp 1666464484
transform 1 0 27324 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_297
timestamp 1666464484
transform 1 0 28428 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_309
timestamp 1666464484
transform 1 0 29532 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_321
timestamp 1666464484
transform 1 0 30636 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_326
timestamp 1666464484
transform 1 0 31096 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_338
timestamp 1666464484
transform 1 0 32200 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_350
timestamp 1666464484
transform 1 0 33304 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_362
timestamp 1666464484
transform 1 0 34408 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_374
timestamp 1666464484
transform 1 0 35512 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_386
timestamp 1666464484
transform 1 0 36616 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_391
timestamp 1666464484
transform 1 0 37076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_403
timestamp 1666464484
transform 1 0 38180 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_415
timestamp 1666464484
transform 1 0 39284 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_427
timestamp 1666464484
transform 1 0 40388 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_439
timestamp 1666464484
transform 1 0 41492 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_451
timestamp 1666464484
transform 1 0 42596 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_456
timestamp 1666464484
transform 1 0 43056 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_468
timestamp 1666464484
transform 1 0 44160 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_480
timestamp 1666464484
transform 1 0 45264 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_492
timestamp 1666464484
transform 1 0 46368 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_504
timestamp 1666464484
transform 1 0 47472 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_516
timestamp 1666464484
transform 1 0 48576 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_521
timestamp 1666464484
transform 1 0 49036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_533
timestamp 1666464484
transform 1 0 50140 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_545
timestamp 1666464484
transform 1 0 51244 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_557
timestamp 1666464484
transform 1 0 52348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_569
timestamp 1666464484
transform 1 0 53452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_581
timestamp 1666464484
transform 1 0 54556 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_586
timestamp 1666464484
transform 1 0 55016 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_598
timestamp 1666464484
transform 1 0 56120 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_610
timestamp 1666464484
transform 1 0 57224 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_622
timestamp 1666464484
transform 1 0 58328 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666464484
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_31
timestamp 1666464484
transform 1 0 3956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_33
timestamp 1666464484
transform 1 0 4140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_45
timestamp 1666464484
transform 1 0 5244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_57
timestamp 1666464484
transform 1 0 6348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_69
timestamp 1666464484
transform 1 0 7452 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_81
timestamp 1666464484
transform 1 0 8556 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_93
timestamp 1666464484
transform 1 0 9660 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_98
timestamp 1666464484
transform 1 0 10120 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_110
timestamp 1666464484
transform 1 0 11224 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_122
timestamp 1666464484
transform 1 0 12328 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_134
timestamp 1666464484
transform 1 0 13432 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_146
timestamp 1666464484
transform 1 0 14536 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_158
timestamp 1666464484
transform 1 0 15640 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_163
timestamp 1666464484
transform 1 0 16100 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_175
timestamp 1666464484
transform 1 0 17204 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_187
timestamp 1666464484
transform 1 0 18308 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_199
timestamp 1666464484
transform 1 0 19412 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_211
timestamp 1666464484
transform 1 0 20516 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_223
timestamp 1666464484
transform 1 0 21620 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_228
timestamp 1666464484
transform 1 0 22080 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_240
timestamp 1666464484
transform 1 0 23184 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_252
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_264
timestamp 1666464484
transform 1 0 25392 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_276
timestamp 1666464484
transform 1 0 26496 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_288
timestamp 1666464484
transform 1 0 27600 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_293
timestamp 1666464484
transform 1 0 28060 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_305
timestamp 1666464484
transform 1 0 29164 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_317
timestamp 1666464484
transform 1 0 30268 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_329
timestamp 1666464484
transform 1 0 31372 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_341
timestamp 1666464484
transform 1 0 32476 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_353
timestamp 1666464484
transform 1 0 33580 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_358
timestamp 1666464484
transform 1 0 34040 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_370
timestamp 1666464484
transform 1 0 35144 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_382
timestamp 1666464484
transform 1 0 36248 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_394
timestamp 1666464484
transform 1 0 37352 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_406
timestamp 1666464484
transform 1 0 38456 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_418
timestamp 1666464484
transform 1 0 39560 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_423
timestamp 1666464484
transform 1 0 40020 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_435
timestamp 1666464484
transform 1 0 41124 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_447
timestamp 1666464484
transform 1 0 42228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_459
timestamp 1666464484
transform 1 0 43332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_471
timestamp 1666464484
transform 1 0 44436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_483
timestamp 1666464484
transform 1 0 45540 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_488
timestamp 1666464484
transform 1 0 46000 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_500
timestamp 1666464484
transform 1 0 47104 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_512
timestamp 1666464484
transform 1 0 48208 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_524
timestamp 1666464484
transform 1 0 49312 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_536
timestamp 1666464484
transform 1 0 50416 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_548
timestamp 1666464484
transform 1 0 51520 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_553
timestamp 1666464484
transform 1 0 51980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_565
timestamp 1666464484
transform 1 0 53084 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_577
timestamp 1666464484
transform 1 0 54188 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1666464484
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1666464484
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_613
timestamp 1666464484
transform 1 0 57500 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_618
timestamp 1666464484
transform 1 0 57960 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_624
timestamp 1666464484
transform 1 0 58512 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666464484
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_51
timestamp 1666464484
transform 1 0 5796 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_63
timestamp 1666464484
transform 1 0 6900 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_66
timestamp 1666464484
transform 1 0 7176 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_78
timestamp 1666464484
transform 1 0 8280 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_90
timestamp 1666464484
transform 1 0 9384 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_102
timestamp 1666464484
transform 1 0 10488 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_114
timestamp 1666464484
transform 1 0 11592 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_126
timestamp 1666464484
transform 1 0 12696 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_131
timestamp 1666464484
transform 1 0 13156 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_143
timestamp 1666464484
transform 1 0 14260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_155
timestamp 1666464484
transform 1 0 15364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_179
timestamp 1666464484
transform 1 0 17572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_191
timestamp 1666464484
transform 1 0 18676 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_196
timestamp 1666464484
transform 1 0 19136 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_208
timestamp 1666464484
transform 1 0 20240 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_220
timestamp 1666464484
transform 1 0 21344 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_232
timestamp 1666464484
transform 1 0 22448 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_244
timestamp 1666464484
transform 1 0 23552 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_256
timestamp 1666464484
transform 1 0 24656 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1666464484
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_273
timestamp 1666464484
transform 1 0 26220 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_285
timestamp 1666464484
transform 1 0 27324 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_297
timestamp 1666464484
transform 1 0 28428 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_309
timestamp 1666464484
transform 1 0 29532 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_321
timestamp 1666464484
transform 1 0 30636 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_326
timestamp 1666464484
transform 1 0 31096 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_338
timestamp 1666464484
transform 1 0 32200 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_350
timestamp 1666464484
transform 1 0 33304 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_362
timestamp 1666464484
transform 1 0 34408 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_374
timestamp 1666464484
transform 1 0 35512 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_386
timestamp 1666464484
transform 1 0 36616 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_391
timestamp 1666464484
transform 1 0 37076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_403
timestamp 1666464484
transform 1 0 38180 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_415
timestamp 1666464484
transform 1 0 39284 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_427
timestamp 1666464484
transform 1 0 40388 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_439
timestamp 1666464484
transform 1 0 41492 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_451
timestamp 1666464484
transform 1 0 42596 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_456
timestamp 1666464484
transform 1 0 43056 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_468
timestamp 1666464484
transform 1 0 44160 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_480
timestamp 1666464484
transform 1 0 45264 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_492
timestamp 1666464484
transform 1 0 46368 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_504
timestamp 1666464484
transform 1 0 47472 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_516
timestamp 1666464484
transform 1 0 48576 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_521
timestamp 1666464484
transform 1 0 49036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_533
timestamp 1666464484
transform 1 0 50140 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_545
timestamp 1666464484
transform 1 0 51244 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_557
timestamp 1666464484
transform 1 0 52348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_569
timestamp 1666464484
transform 1 0 53452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_581
timestamp 1666464484
transform 1 0 54556 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_586
timestamp 1666464484
transform 1 0 55016 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_598
timestamp 1666464484
transform 1 0 56120 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_610
timestamp 1666464484
transform 1 0 57224 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_622
timestamp 1666464484
transform 1 0 58328 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666464484
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1666464484
transform 1 0 3588 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_31
timestamp 1666464484
transform 1 0 3956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_33
timestamp 1666464484
transform 1 0 4140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_45
timestamp 1666464484
transform 1 0 5244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_57
timestamp 1666464484
transform 1 0 6348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_69
timestamp 1666464484
transform 1 0 7452 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_81
timestamp 1666464484
transform 1 0 8556 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_93
timestamp 1666464484
transform 1 0 9660 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_98
timestamp 1666464484
transform 1 0 10120 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_110
timestamp 1666464484
transform 1 0 11224 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_122
timestamp 1666464484
transform 1 0 12328 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_134
timestamp 1666464484
transform 1 0 13432 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_146
timestamp 1666464484
transform 1 0 14536 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_158
timestamp 1666464484
transform 1 0 15640 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_163
timestamp 1666464484
transform 1 0 16100 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_175
timestamp 1666464484
transform 1 0 17204 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_187
timestamp 1666464484
transform 1 0 18308 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_199
timestamp 1666464484
transform 1 0 19412 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_211
timestamp 1666464484
transform 1 0 20516 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_223
timestamp 1666464484
transform 1 0 21620 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_228
timestamp 1666464484
transform 1 0 22080 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_240
timestamp 1666464484
transform 1 0 23184 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_252
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_264
timestamp 1666464484
transform 1 0 25392 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_276
timestamp 1666464484
transform 1 0 26496 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_288
timestamp 1666464484
transform 1 0 27600 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_293
timestamp 1666464484
transform 1 0 28060 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_305
timestamp 1666464484
transform 1 0 29164 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_317
timestamp 1666464484
transform 1 0 30268 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_329
timestamp 1666464484
transform 1 0 31372 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_341
timestamp 1666464484
transform 1 0 32476 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_353
timestamp 1666464484
transform 1 0 33580 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_358
timestamp 1666464484
transform 1 0 34040 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_370
timestamp 1666464484
transform 1 0 35144 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_382
timestamp 1666464484
transform 1 0 36248 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_394
timestamp 1666464484
transform 1 0 37352 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_406
timestamp 1666464484
transform 1 0 38456 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_418
timestamp 1666464484
transform 1 0 39560 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_423
timestamp 1666464484
transform 1 0 40020 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_435
timestamp 1666464484
transform 1 0 41124 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_447
timestamp 1666464484
transform 1 0 42228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_459
timestamp 1666464484
transform 1 0 43332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_471
timestamp 1666464484
transform 1 0 44436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_483
timestamp 1666464484
transform 1 0 45540 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_488
timestamp 1666464484
transform 1 0 46000 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_500
timestamp 1666464484
transform 1 0 47104 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_512
timestamp 1666464484
transform 1 0 48208 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_524
timestamp 1666464484
transform 1 0 49312 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_536
timestamp 1666464484
transform 1 0 50416 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_548
timestamp 1666464484
transform 1 0 51520 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_553
timestamp 1666464484
transform 1 0 51980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_565
timestamp 1666464484
transform 1 0 53084 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_577
timestamp 1666464484
transform 1 0 54188 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1666464484
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1666464484
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_613
timestamp 1666464484
transform 1 0 57500 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_618
timestamp 1666464484
transform 1 0 57960 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_624
timestamp 1666464484
transform 1 0 58512 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666464484
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1666464484
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1666464484
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_51
timestamp 1666464484
transform 1 0 5796 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_63
timestamp 1666464484
transform 1 0 6900 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_66
timestamp 1666464484
transform 1 0 7176 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_78
timestamp 1666464484
transform 1 0 8280 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_90
timestamp 1666464484
transform 1 0 9384 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_102
timestamp 1666464484
transform 1 0 10488 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_114
timestamp 1666464484
transform 1 0 11592 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_126
timestamp 1666464484
transform 1 0 12696 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_131
timestamp 1666464484
transform 1 0 13156 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_143
timestamp 1666464484
transform 1 0 14260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_155
timestamp 1666464484
transform 1 0 15364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_167
timestamp 1666464484
transform 1 0 16468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_179
timestamp 1666464484
transform 1 0 17572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_191
timestamp 1666464484
transform 1 0 18676 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_196
timestamp 1666464484
transform 1 0 19136 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_208
timestamp 1666464484
transform 1 0 20240 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_220
timestamp 1666464484
transform 1 0 21344 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_232
timestamp 1666464484
transform 1 0 22448 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_244
timestamp 1666464484
transform 1 0 23552 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_256
timestamp 1666464484
transform 1 0 24656 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1666464484
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_273
timestamp 1666464484
transform 1 0 26220 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_285
timestamp 1666464484
transform 1 0 27324 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_297
timestamp 1666464484
transform 1 0 28428 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_309
timestamp 1666464484
transform 1 0 29532 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_321
timestamp 1666464484
transform 1 0 30636 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_326
timestamp 1666464484
transform 1 0 31096 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_338
timestamp 1666464484
transform 1 0 32200 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_350
timestamp 1666464484
transform 1 0 33304 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_362
timestamp 1666464484
transform 1 0 34408 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_374
timestamp 1666464484
transform 1 0 35512 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_386
timestamp 1666464484
transform 1 0 36616 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_391
timestamp 1666464484
transform 1 0 37076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_403
timestamp 1666464484
transform 1 0 38180 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_415
timestamp 1666464484
transform 1 0 39284 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_427
timestamp 1666464484
transform 1 0 40388 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_439
timestamp 1666464484
transform 1 0 41492 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_451
timestamp 1666464484
transform 1 0 42596 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_456
timestamp 1666464484
transform 1 0 43056 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_468
timestamp 1666464484
transform 1 0 44160 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_480
timestamp 1666464484
transform 1 0 45264 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_492
timestamp 1666464484
transform 1 0 46368 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_504
timestamp 1666464484
transform 1 0 47472 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_516
timestamp 1666464484
transform 1 0 48576 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_521
timestamp 1666464484
transform 1 0 49036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_533
timestamp 1666464484
transform 1 0 50140 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_545
timestamp 1666464484
transform 1 0 51244 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_557
timestamp 1666464484
transform 1 0 52348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_569
timestamp 1666464484
transform 1 0 53452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_581
timestamp 1666464484
transform 1 0 54556 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_586
timestamp 1666464484
transform 1 0 55016 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_598
timestamp 1666464484
transform 1 0 56120 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_610
timestamp 1666464484
transform 1 0 57224 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_622
timestamp 1666464484
transform 1 0 58328 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1666464484
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1666464484
transform 1 0 3588 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_31
timestamp 1666464484
transform 1 0 3956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_33
timestamp 1666464484
transform 1 0 4140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_45
timestamp 1666464484
transform 1 0 5244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_57
timestamp 1666464484
transform 1 0 6348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_69
timestamp 1666464484
transform 1 0 7452 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_81
timestamp 1666464484
transform 1 0 8556 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_93
timestamp 1666464484
transform 1 0 9660 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_98
timestamp 1666464484
transform 1 0 10120 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_110
timestamp 1666464484
transform 1 0 11224 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_122
timestamp 1666464484
transform 1 0 12328 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_134
timestamp 1666464484
transform 1 0 13432 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_146
timestamp 1666464484
transform 1 0 14536 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_158
timestamp 1666464484
transform 1 0 15640 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_163
timestamp 1666464484
transform 1 0 16100 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_175
timestamp 1666464484
transform 1 0 17204 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_187
timestamp 1666464484
transform 1 0 18308 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_199
timestamp 1666464484
transform 1 0 19412 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_211
timestamp 1666464484
transform 1 0 20516 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_223
timestamp 1666464484
transform 1 0 21620 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_228
timestamp 1666464484
transform 1 0 22080 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_240
timestamp 1666464484
transform 1 0 23184 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_252
timestamp 1666464484
transform 1 0 24288 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_264
timestamp 1666464484
transform 1 0 25392 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_276
timestamp 1666464484
transform 1 0 26496 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_288
timestamp 1666464484
transform 1 0 27600 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_293
timestamp 1666464484
transform 1 0 28060 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_305
timestamp 1666464484
transform 1 0 29164 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_317
timestamp 1666464484
transform 1 0 30268 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_329
timestamp 1666464484
transform 1 0 31372 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_341
timestamp 1666464484
transform 1 0 32476 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_353
timestamp 1666464484
transform 1 0 33580 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_358
timestamp 1666464484
transform 1 0 34040 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_370
timestamp 1666464484
transform 1 0 35144 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_382
timestamp 1666464484
transform 1 0 36248 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_394
timestamp 1666464484
transform 1 0 37352 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_406
timestamp 1666464484
transform 1 0 38456 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_418
timestamp 1666464484
transform 1 0 39560 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_423
timestamp 1666464484
transform 1 0 40020 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_435
timestamp 1666464484
transform 1 0 41124 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_447
timestamp 1666464484
transform 1 0 42228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_459
timestamp 1666464484
transform 1 0 43332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_471
timestamp 1666464484
transform 1 0 44436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_483
timestamp 1666464484
transform 1 0 45540 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_488
timestamp 1666464484
transform 1 0 46000 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_500
timestamp 1666464484
transform 1 0 47104 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_512
timestamp 1666464484
transform 1 0 48208 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_524
timestamp 1666464484
transform 1 0 49312 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_536
timestamp 1666464484
transform 1 0 50416 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_548
timestamp 1666464484
transform 1 0 51520 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_553
timestamp 1666464484
transform 1 0 51980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_565
timestamp 1666464484
transform 1 0 53084 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_577
timestamp 1666464484
transform 1 0 54188 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1666464484
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1666464484
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_613
timestamp 1666464484
transform 1 0 57500 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_618
timestamp 1666464484
transform 1 0 57960 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_624
timestamp 1666464484
transform 1 0 58512 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666464484
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666464484
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1666464484
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_51
timestamp 1666464484
transform 1 0 5796 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_63
timestamp 1666464484
transform 1 0 6900 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_66
timestamp 1666464484
transform 1 0 7176 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_78
timestamp 1666464484
transform 1 0 8280 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_90
timestamp 1666464484
transform 1 0 9384 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_102
timestamp 1666464484
transform 1 0 10488 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_114
timestamp 1666464484
transform 1 0 11592 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_126
timestamp 1666464484
transform 1 0 12696 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_131
timestamp 1666464484
transform 1 0 13156 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_143
timestamp 1666464484
transform 1 0 14260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_155
timestamp 1666464484
transform 1 0 15364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_167
timestamp 1666464484
transform 1 0 16468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_179
timestamp 1666464484
transform 1 0 17572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_191
timestamp 1666464484
transform 1 0 18676 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_196
timestamp 1666464484
transform 1 0 19136 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_208
timestamp 1666464484
transform 1 0 20240 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_220
timestamp 1666464484
transform 1 0 21344 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_232
timestamp 1666464484
transform 1 0 22448 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_244
timestamp 1666464484
transform 1 0 23552 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_256
timestamp 1666464484
transform 1 0 24656 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1666464484
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_273
timestamp 1666464484
transform 1 0 26220 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_285
timestamp 1666464484
transform 1 0 27324 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_297
timestamp 1666464484
transform 1 0 28428 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_309
timestamp 1666464484
transform 1 0 29532 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_321
timestamp 1666464484
transform 1 0 30636 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_326
timestamp 1666464484
transform 1 0 31096 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_338
timestamp 1666464484
transform 1 0 32200 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_350
timestamp 1666464484
transform 1 0 33304 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_362
timestamp 1666464484
transform 1 0 34408 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_374
timestamp 1666464484
transform 1 0 35512 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_386
timestamp 1666464484
transform 1 0 36616 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_391
timestamp 1666464484
transform 1 0 37076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_403
timestamp 1666464484
transform 1 0 38180 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_415
timestamp 1666464484
transform 1 0 39284 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_427
timestamp 1666464484
transform 1 0 40388 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_439
timestamp 1666464484
transform 1 0 41492 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_451
timestamp 1666464484
transform 1 0 42596 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_456
timestamp 1666464484
transform 1 0 43056 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_468
timestamp 1666464484
transform 1 0 44160 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_480
timestamp 1666464484
transform 1 0 45264 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_492
timestamp 1666464484
transform 1 0 46368 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_504
timestamp 1666464484
transform 1 0 47472 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_516
timestamp 1666464484
transform 1 0 48576 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_521
timestamp 1666464484
transform 1 0 49036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_533
timestamp 1666464484
transform 1 0 50140 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_545
timestamp 1666464484
transform 1 0 51244 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_557
timestamp 1666464484
transform 1 0 52348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_569
timestamp 1666464484
transform 1 0 53452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_581
timestamp 1666464484
transform 1 0 54556 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_586
timestamp 1666464484
transform 1 0 55016 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_598
timestamp 1666464484
transform 1 0 56120 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_610
timestamp 1666464484
transform 1 0 57224 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_622
timestamp 1666464484
transform 1 0 58328 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1666464484
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1666464484
transform 1 0 3588 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_31
timestamp 1666464484
transform 1 0 3956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_33
timestamp 1666464484
transform 1 0 4140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_45
timestamp 1666464484
transform 1 0 5244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_57
timestamp 1666464484
transform 1 0 6348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_69
timestamp 1666464484
transform 1 0 7452 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_81
timestamp 1666464484
transform 1 0 8556 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_93
timestamp 1666464484
transform 1 0 9660 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_98
timestamp 1666464484
transform 1 0 10120 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_110
timestamp 1666464484
transform 1 0 11224 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_122
timestamp 1666464484
transform 1 0 12328 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_134
timestamp 1666464484
transform 1 0 13432 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_146
timestamp 1666464484
transform 1 0 14536 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_158
timestamp 1666464484
transform 1 0 15640 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_163
timestamp 1666464484
transform 1 0 16100 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_175
timestamp 1666464484
transform 1 0 17204 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_187
timestamp 1666464484
transform 1 0 18308 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_199
timestamp 1666464484
transform 1 0 19412 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_211
timestamp 1666464484
transform 1 0 20516 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_223
timestamp 1666464484
transform 1 0 21620 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_228
timestamp 1666464484
transform 1 0 22080 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_240
timestamp 1666464484
transform 1 0 23184 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_252
timestamp 1666464484
transform 1 0 24288 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_264
timestamp 1666464484
transform 1 0 25392 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_276
timestamp 1666464484
transform 1 0 26496 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_288
timestamp 1666464484
transform 1 0 27600 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_293
timestamp 1666464484
transform 1 0 28060 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_305
timestamp 1666464484
transform 1 0 29164 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_317
timestamp 1666464484
transform 1 0 30268 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_329
timestamp 1666464484
transform 1 0 31372 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_341
timestamp 1666464484
transform 1 0 32476 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_353
timestamp 1666464484
transform 1 0 33580 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_358
timestamp 1666464484
transform 1 0 34040 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_370
timestamp 1666464484
transform 1 0 35144 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_382
timestamp 1666464484
transform 1 0 36248 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_394
timestamp 1666464484
transform 1 0 37352 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_406
timestamp 1666464484
transform 1 0 38456 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_418
timestamp 1666464484
transform 1 0 39560 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_423
timestamp 1666464484
transform 1 0 40020 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_435
timestamp 1666464484
transform 1 0 41124 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_447
timestamp 1666464484
transform 1 0 42228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_459
timestamp 1666464484
transform 1 0 43332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_471
timestamp 1666464484
transform 1 0 44436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_483
timestamp 1666464484
transform 1 0 45540 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_488
timestamp 1666464484
transform 1 0 46000 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_500
timestamp 1666464484
transform 1 0 47104 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_512
timestamp 1666464484
transform 1 0 48208 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_524
timestamp 1666464484
transform 1 0 49312 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_536
timestamp 1666464484
transform 1 0 50416 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_548
timestamp 1666464484
transform 1 0 51520 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_553
timestamp 1666464484
transform 1 0 51980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_565
timestamp 1666464484
transform 1 0 53084 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_577
timestamp 1666464484
transform 1 0 54188 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1666464484
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1666464484
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_613
timestamp 1666464484
transform 1 0 57500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_618
timestamp 1666464484
transform 1 0 57960 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_624
timestamp 1666464484
transform 1 0 58512 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666464484
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1666464484
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1666464484
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_51
timestamp 1666464484
transform 1 0 5796 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_63
timestamp 1666464484
transform 1 0 6900 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_66
timestamp 1666464484
transform 1 0 7176 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_78
timestamp 1666464484
transform 1 0 8280 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_90
timestamp 1666464484
transform 1 0 9384 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_102
timestamp 1666464484
transform 1 0 10488 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_114
timestamp 1666464484
transform 1 0 11592 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_126
timestamp 1666464484
transform 1 0 12696 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_131
timestamp 1666464484
transform 1 0 13156 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_143
timestamp 1666464484
transform 1 0 14260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_155
timestamp 1666464484
transform 1 0 15364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_167
timestamp 1666464484
transform 1 0 16468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_179
timestamp 1666464484
transform 1 0 17572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_191
timestamp 1666464484
transform 1 0 18676 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_196
timestamp 1666464484
transform 1 0 19136 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_208
timestamp 1666464484
transform 1 0 20240 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_220
timestamp 1666464484
transform 1 0 21344 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_232
timestamp 1666464484
transform 1 0 22448 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_244
timestamp 1666464484
transform 1 0 23552 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_256
timestamp 1666464484
transform 1 0 24656 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1666464484
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_273
timestamp 1666464484
transform 1 0 26220 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_285
timestamp 1666464484
transform 1 0 27324 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_297
timestamp 1666464484
transform 1 0 28428 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_309
timestamp 1666464484
transform 1 0 29532 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_321
timestamp 1666464484
transform 1 0 30636 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_326
timestamp 1666464484
transform 1 0 31096 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_338
timestamp 1666464484
transform 1 0 32200 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_350
timestamp 1666464484
transform 1 0 33304 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_362
timestamp 1666464484
transform 1 0 34408 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_374
timestamp 1666464484
transform 1 0 35512 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_386
timestamp 1666464484
transform 1 0 36616 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_391
timestamp 1666464484
transform 1 0 37076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_403
timestamp 1666464484
transform 1 0 38180 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_415
timestamp 1666464484
transform 1 0 39284 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_427
timestamp 1666464484
transform 1 0 40388 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_439
timestamp 1666464484
transform 1 0 41492 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_451
timestamp 1666464484
transform 1 0 42596 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_456
timestamp 1666464484
transform 1 0 43056 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_468
timestamp 1666464484
transform 1 0 44160 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_480
timestamp 1666464484
transform 1 0 45264 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_492
timestamp 1666464484
transform 1 0 46368 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_504
timestamp 1666464484
transform 1 0 47472 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_516
timestamp 1666464484
transform 1 0 48576 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_521
timestamp 1666464484
transform 1 0 49036 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_533
timestamp 1666464484
transform 1 0 50140 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_545
timestamp 1666464484
transform 1 0 51244 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_557
timestamp 1666464484
transform 1 0 52348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_569
timestamp 1666464484
transform 1 0 53452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_581
timestamp 1666464484
transform 1 0 54556 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_586
timestamp 1666464484
transform 1 0 55016 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_598
timestamp 1666464484
transform 1 0 56120 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_610
timestamp 1666464484
transform 1 0 57224 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_622
timestamp 1666464484
transform 1 0 58328 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1666464484
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1666464484
transform 1 0 3588 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_31
timestamp 1666464484
transform 1 0 3956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_33
timestamp 1666464484
transform 1 0 4140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_45
timestamp 1666464484
transform 1 0 5244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_57
timestamp 1666464484
transform 1 0 6348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_69
timestamp 1666464484
transform 1 0 7452 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_81
timestamp 1666464484
transform 1 0 8556 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_93
timestamp 1666464484
transform 1 0 9660 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_98
timestamp 1666464484
transform 1 0 10120 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_110
timestamp 1666464484
transform 1 0 11224 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_122
timestamp 1666464484
transform 1 0 12328 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_134
timestamp 1666464484
transform 1 0 13432 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_146
timestamp 1666464484
transform 1 0 14536 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_158
timestamp 1666464484
transform 1 0 15640 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_163
timestamp 1666464484
transform 1 0 16100 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_175
timestamp 1666464484
transform 1 0 17204 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_187
timestamp 1666464484
transform 1 0 18308 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_199
timestamp 1666464484
transform 1 0 19412 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_211
timestamp 1666464484
transform 1 0 20516 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_223
timestamp 1666464484
transform 1 0 21620 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_228
timestamp 1666464484
transform 1 0 22080 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_240
timestamp 1666464484
transform 1 0 23184 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_252
timestamp 1666464484
transform 1 0 24288 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_264
timestamp 1666464484
transform 1 0 25392 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_276
timestamp 1666464484
transform 1 0 26496 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_288
timestamp 1666464484
transform 1 0 27600 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_293
timestamp 1666464484
transform 1 0 28060 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_305
timestamp 1666464484
transform 1 0 29164 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_317
timestamp 1666464484
transform 1 0 30268 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_329
timestamp 1666464484
transform 1 0 31372 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_341
timestamp 1666464484
transform 1 0 32476 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_353
timestamp 1666464484
transform 1 0 33580 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_358
timestamp 1666464484
transform 1 0 34040 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_370
timestamp 1666464484
transform 1 0 35144 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_382
timestamp 1666464484
transform 1 0 36248 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_394
timestamp 1666464484
transform 1 0 37352 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_406
timestamp 1666464484
transform 1 0 38456 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_418
timestamp 1666464484
transform 1 0 39560 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_423
timestamp 1666464484
transform 1 0 40020 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_435
timestamp 1666464484
transform 1 0 41124 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_447
timestamp 1666464484
transform 1 0 42228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_459
timestamp 1666464484
transform 1 0 43332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_471
timestamp 1666464484
transform 1 0 44436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_483
timestamp 1666464484
transform 1 0 45540 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_488
timestamp 1666464484
transform 1 0 46000 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_500
timestamp 1666464484
transform 1 0 47104 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_512
timestamp 1666464484
transform 1 0 48208 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_524
timestamp 1666464484
transform 1 0 49312 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_536
timestamp 1666464484
transform 1 0 50416 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_548
timestamp 1666464484
transform 1 0 51520 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_553
timestamp 1666464484
transform 1 0 51980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_565
timestamp 1666464484
transform 1 0 53084 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_577
timestamp 1666464484
transform 1 0 54188 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1666464484
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1666464484
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_613
timestamp 1666464484
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_618
timestamp 1666464484
transform 1 0 57960 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_624
timestamp 1666464484
transform 1 0 58512 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666464484
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1666464484
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1666464484
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_51
timestamp 1666464484
transform 1 0 5796 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_63
timestamp 1666464484
transform 1 0 6900 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_66
timestamp 1666464484
transform 1 0 7176 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_78
timestamp 1666464484
transform 1 0 8280 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_90
timestamp 1666464484
transform 1 0 9384 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_102
timestamp 1666464484
transform 1 0 10488 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_114
timestamp 1666464484
transform 1 0 11592 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_126
timestamp 1666464484
transform 1 0 12696 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_131
timestamp 1666464484
transform 1 0 13156 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_143
timestamp 1666464484
transform 1 0 14260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_155
timestamp 1666464484
transform 1 0 15364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_167
timestamp 1666464484
transform 1 0 16468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_179
timestamp 1666464484
transform 1 0 17572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_191
timestamp 1666464484
transform 1 0 18676 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_196
timestamp 1666464484
transform 1 0 19136 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_208
timestamp 1666464484
transform 1 0 20240 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_220
timestamp 1666464484
transform 1 0 21344 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_232
timestamp 1666464484
transform 1 0 22448 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_244
timestamp 1666464484
transform 1 0 23552 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_256
timestamp 1666464484
transform 1 0 24656 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1666464484
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_273
timestamp 1666464484
transform 1 0 26220 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_285
timestamp 1666464484
transform 1 0 27324 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_297
timestamp 1666464484
transform 1 0 28428 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_309
timestamp 1666464484
transform 1 0 29532 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_321
timestamp 1666464484
transform 1 0 30636 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_326
timestamp 1666464484
transform 1 0 31096 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_338
timestamp 1666464484
transform 1 0 32200 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_350
timestamp 1666464484
transform 1 0 33304 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_362
timestamp 1666464484
transform 1 0 34408 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_374
timestamp 1666464484
transform 1 0 35512 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_386
timestamp 1666464484
transform 1 0 36616 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_391
timestamp 1666464484
transform 1 0 37076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_403
timestamp 1666464484
transform 1 0 38180 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_415
timestamp 1666464484
transform 1 0 39284 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_427
timestamp 1666464484
transform 1 0 40388 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_439
timestamp 1666464484
transform 1 0 41492 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_451
timestamp 1666464484
transform 1 0 42596 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_456
timestamp 1666464484
transform 1 0 43056 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_468
timestamp 1666464484
transform 1 0 44160 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_480
timestamp 1666464484
transform 1 0 45264 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_492
timestamp 1666464484
transform 1 0 46368 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_504
timestamp 1666464484
transform 1 0 47472 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_516
timestamp 1666464484
transform 1 0 48576 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_521
timestamp 1666464484
transform 1 0 49036 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_533
timestamp 1666464484
transform 1 0 50140 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_545
timestamp 1666464484
transform 1 0 51244 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_557
timestamp 1666464484
transform 1 0 52348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_569
timestamp 1666464484
transform 1 0 53452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_581
timestamp 1666464484
transform 1 0 54556 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_586
timestamp 1666464484
transform 1 0 55016 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_598
timestamp 1666464484
transform 1 0 56120 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_610
timestamp 1666464484
transform 1 0 57224 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_622
timestamp 1666464484
transform 1 0 58328 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1666464484
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1666464484
transform 1 0 3588 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_31
timestamp 1666464484
transform 1 0 3956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_33
timestamp 1666464484
transform 1 0 4140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_45
timestamp 1666464484
transform 1 0 5244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_57
timestamp 1666464484
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_69
timestamp 1666464484
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_81
timestamp 1666464484
transform 1 0 8556 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_93
timestamp 1666464484
transform 1 0 9660 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_98
timestamp 1666464484
transform 1 0 10120 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_110
timestamp 1666464484
transform 1 0 11224 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_122
timestamp 1666464484
transform 1 0 12328 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_134
timestamp 1666464484
transform 1 0 13432 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_146
timestamp 1666464484
transform 1 0 14536 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_158
timestamp 1666464484
transform 1 0 15640 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_163
timestamp 1666464484
transform 1 0 16100 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_175
timestamp 1666464484
transform 1 0 17204 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_187
timestamp 1666464484
transform 1 0 18308 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_199
timestamp 1666464484
transform 1 0 19412 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_211
timestamp 1666464484
transform 1 0 20516 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_223
timestamp 1666464484
transform 1 0 21620 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_228
timestamp 1666464484
transform 1 0 22080 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_240
timestamp 1666464484
transform 1 0 23184 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_252
timestamp 1666464484
transform 1 0 24288 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_264
timestamp 1666464484
transform 1 0 25392 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_276
timestamp 1666464484
transform 1 0 26496 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_288
timestamp 1666464484
transform 1 0 27600 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_293
timestamp 1666464484
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_305
timestamp 1666464484
transform 1 0 29164 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_317
timestamp 1666464484
transform 1 0 30268 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_329
timestamp 1666464484
transform 1 0 31372 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_341
timestamp 1666464484
transform 1 0 32476 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_353
timestamp 1666464484
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_358
timestamp 1666464484
transform 1 0 34040 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_370
timestamp 1666464484
transform 1 0 35144 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_382
timestamp 1666464484
transform 1 0 36248 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_394
timestamp 1666464484
transform 1 0 37352 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_406
timestamp 1666464484
transform 1 0 38456 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_418
timestamp 1666464484
transform 1 0 39560 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_423
timestamp 1666464484
transform 1 0 40020 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_435
timestamp 1666464484
transform 1 0 41124 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_447
timestamp 1666464484
transform 1 0 42228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_459
timestamp 1666464484
transform 1 0 43332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_471
timestamp 1666464484
transform 1 0 44436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_483
timestamp 1666464484
transform 1 0 45540 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_488
timestamp 1666464484
transform 1 0 46000 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_500
timestamp 1666464484
transform 1 0 47104 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_512
timestamp 1666464484
transform 1 0 48208 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_524
timestamp 1666464484
transform 1 0 49312 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_536
timestamp 1666464484
transform 1 0 50416 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_548
timestamp 1666464484
transform 1 0 51520 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_553
timestamp 1666464484
transform 1 0 51980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_565
timestamp 1666464484
transform 1 0 53084 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_577
timestamp 1666464484
transform 1 0 54188 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1666464484
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1666464484
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_613
timestamp 1666464484
transform 1 0 57500 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_618
timestamp 1666464484
transform 1 0 57960 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_624
timestamp 1666464484
transform 1 0 58512 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1666464484
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1666464484
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1666464484
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1666464484
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_51
timestamp 1666464484
transform 1 0 5796 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_63
timestamp 1666464484
transform 1 0 6900 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_66
timestamp 1666464484
transform 1 0 7176 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_78
timestamp 1666464484
transform 1 0 8280 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_90
timestamp 1666464484
transform 1 0 9384 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_102
timestamp 1666464484
transform 1 0 10488 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_114
timestamp 1666464484
transform 1 0 11592 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_126
timestamp 1666464484
transform 1 0 12696 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_131
timestamp 1666464484
transform 1 0 13156 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_143
timestamp 1666464484
transform 1 0 14260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_155
timestamp 1666464484
transform 1 0 15364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_167
timestamp 1666464484
transform 1 0 16468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_179
timestamp 1666464484
transform 1 0 17572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_191
timestamp 1666464484
transform 1 0 18676 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_196
timestamp 1666464484
transform 1 0 19136 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_208
timestamp 1666464484
transform 1 0 20240 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_220
timestamp 1666464484
transform 1 0 21344 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_232
timestamp 1666464484
transform 1 0 22448 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_244
timestamp 1666464484
transform 1 0 23552 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_256
timestamp 1666464484
transform 1 0 24656 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1666464484
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_273
timestamp 1666464484
transform 1 0 26220 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_285
timestamp 1666464484
transform 1 0 27324 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_297
timestamp 1666464484
transform 1 0 28428 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_309
timestamp 1666464484
transform 1 0 29532 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_321
timestamp 1666464484
transform 1 0 30636 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_326
timestamp 1666464484
transform 1 0 31096 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_338
timestamp 1666464484
transform 1 0 32200 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_350
timestamp 1666464484
transform 1 0 33304 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_362
timestamp 1666464484
transform 1 0 34408 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_374
timestamp 1666464484
transform 1 0 35512 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_386
timestamp 1666464484
transform 1 0 36616 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_391
timestamp 1666464484
transform 1 0 37076 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_403
timestamp 1666464484
transform 1 0 38180 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_415
timestamp 1666464484
transform 1 0 39284 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_427
timestamp 1666464484
transform 1 0 40388 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_439
timestamp 1666464484
transform 1 0 41492 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_451
timestamp 1666464484
transform 1 0 42596 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_456
timestamp 1666464484
transform 1 0 43056 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_468
timestamp 1666464484
transform 1 0 44160 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_480
timestamp 1666464484
transform 1 0 45264 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_492
timestamp 1666464484
transform 1 0 46368 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_504
timestamp 1666464484
transform 1 0 47472 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_516
timestamp 1666464484
transform 1 0 48576 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_521
timestamp 1666464484
transform 1 0 49036 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_533
timestamp 1666464484
transform 1 0 50140 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_545
timestamp 1666464484
transform 1 0 51244 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_557
timestamp 1666464484
transform 1 0 52348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_569
timestamp 1666464484
transform 1 0 53452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_581
timestamp 1666464484
transform 1 0 54556 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_586
timestamp 1666464484
transform 1 0 55016 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_598
timestamp 1666464484
transform 1 0 56120 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_610
timestamp 1666464484
transform 1 0 57224 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_622
timestamp 1666464484
transform 1 0 58328 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1666464484
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1666464484
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_27
timestamp 1666464484
transform 1 0 3588 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_31
timestamp 1666464484
transform 1 0 3956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_33
timestamp 1666464484
transform 1 0 4140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_45
timestamp 1666464484
transform 1 0 5244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_57
timestamp 1666464484
transform 1 0 6348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_69
timestamp 1666464484
transform 1 0 7452 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_81
timestamp 1666464484
transform 1 0 8556 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_93
timestamp 1666464484
transform 1 0 9660 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_98
timestamp 1666464484
transform 1 0 10120 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_110
timestamp 1666464484
transform 1 0 11224 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_122
timestamp 1666464484
transform 1 0 12328 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_134
timestamp 1666464484
transform 1 0 13432 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_146
timestamp 1666464484
transform 1 0 14536 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_158
timestamp 1666464484
transform 1 0 15640 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_163
timestamp 1666464484
transform 1 0 16100 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_175
timestamp 1666464484
transform 1 0 17204 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_187
timestamp 1666464484
transform 1 0 18308 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_199
timestamp 1666464484
transform 1 0 19412 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_211
timestamp 1666464484
transform 1 0 20516 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_223
timestamp 1666464484
transform 1 0 21620 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_228
timestamp 1666464484
transform 1 0 22080 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_240
timestamp 1666464484
transform 1 0 23184 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_252
timestamp 1666464484
transform 1 0 24288 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_264
timestamp 1666464484
transform 1 0 25392 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_276
timestamp 1666464484
transform 1 0 26496 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_288
timestamp 1666464484
transform 1 0 27600 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_293
timestamp 1666464484
transform 1 0 28060 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_305
timestamp 1666464484
transform 1 0 29164 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_317
timestamp 1666464484
transform 1 0 30268 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_329
timestamp 1666464484
transform 1 0 31372 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_341
timestamp 1666464484
transform 1 0 32476 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_353
timestamp 1666464484
transform 1 0 33580 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_358
timestamp 1666464484
transform 1 0 34040 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_370
timestamp 1666464484
transform 1 0 35144 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_382
timestamp 1666464484
transform 1 0 36248 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_394
timestamp 1666464484
transform 1 0 37352 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_406
timestamp 1666464484
transform 1 0 38456 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_418
timestamp 1666464484
transform 1 0 39560 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_423
timestamp 1666464484
transform 1 0 40020 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_435
timestamp 1666464484
transform 1 0 41124 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_447
timestamp 1666464484
transform 1 0 42228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_459
timestamp 1666464484
transform 1 0 43332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_471
timestamp 1666464484
transform 1 0 44436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_483
timestamp 1666464484
transform 1 0 45540 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_488
timestamp 1666464484
transform 1 0 46000 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_500
timestamp 1666464484
transform 1 0 47104 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_512
timestamp 1666464484
transform 1 0 48208 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_524
timestamp 1666464484
transform 1 0 49312 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_536
timestamp 1666464484
transform 1 0 50416 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_548
timestamp 1666464484
transform 1 0 51520 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_553
timestamp 1666464484
transform 1 0 51980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_565
timestamp 1666464484
transform 1 0 53084 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_577
timestamp 1666464484
transform 1 0 54188 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1666464484
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1666464484
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_613
timestamp 1666464484
transform 1 0 57500 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_618
timestamp 1666464484
transform 1 0 57960 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_624
timestamp 1666464484
transform 1 0 58512 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1666464484
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1666464484
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1666464484
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1666464484
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_51
timestamp 1666464484
transform 1 0 5796 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_63
timestamp 1666464484
transform 1 0 6900 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_66
timestamp 1666464484
transform 1 0 7176 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_78
timestamp 1666464484
transform 1 0 8280 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_90
timestamp 1666464484
transform 1 0 9384 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_102
timestamp 1666464484
transform 1 0 10488 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_114
timestamp 1666464484
transform 1 0 11592 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_126
timestamp 1666464484
transform 1 0 12696 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_131
timestamp 1666464484
transform 1 0 13156 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_143
timestamp 1666464484
transform 1 0 14260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_155
timestamp 1666464484
transform 1 0 15364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_167
timestamp 1666464484
transform 1 0 16468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_179
timestamp 1666464484
transform 1 0 17572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_191
timestamp 1666464484
transform 1 0 18676 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_196
timestamp 1666464484
transform 1 0 19136 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_208
timestamp 1666464484
transform 1 0 20240 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_220
timestamp 1666464484
transform 1 0 21344 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_232
timestamp 1666464484
transform 1 0 22448 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_244
timestamp 1666464484
transform 1 0 23552 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_256
timestamp 1666464484
transform 1 0 24656 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1666464484
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_273
timestamp 1666464484
transform 1 0 26220 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_285
timestamp 1666464484
transform 1 0 27324 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_297
timestamp 1666464484
transform 1 0 28428 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_309
timestamp 1666464484
transform 1 0 29532 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_321
timestamp 1666464484
transform 1 0 30636 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_326
timestamp 1666464484
transform 1 0 31096 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_338
timestamp 1666464484
transform 1 0 32200 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_350
timestamp 1666464484
transform 1 0 33304 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_362
timestamp 1666464484
transform 1 0 34408 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_374
timestamp 1666464484
transform 1 0 35512 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_386
timestamp 1666464484
transform 1 0 36616 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_391
timestamp 1666464484
transform 1 0 37076 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_403
timestamp 1666464484
transform 1 0 38180 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_415
timestamp 1666464484
transform 1 0 39284 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_427
timestamp 1666464484
transform 1 0 40388 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_439
timestamp 1666464484
transform 1 0 41492 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_451
timestamp 1666464484
transform 1 0 42596 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_456
timestamp 1666464484
transform 1 0 43056 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_468
timestamp 1666464484
transform 1 0 44160 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_480
timestamp 1666464484
transform 1 0 45264 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_492
timestamp 1666464484
transform 1 0 46368 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_504
timestamp 1666464484
transform 1 0 47472 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_516
timestamp 1666464484
transform 1 0 48576 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_521
timestamp 1666464484
transform 1 0 49036 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_533
timestamp 1666464484
transform 1 0 50140 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_545
timestamp 1666464484
transform 1 0 51244 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_557
timestamp 1666464484
transform 1 0 52348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_569
timestamp 1666464484
transform 1 0 53452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_581
timestamp 1666464484
transform 1 0 54556 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_586
timestamp 1666464484
transform 1 0 55016 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_598
timestamp 1666464484
transform 1 0 56120 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_610
timestamp 1666464484
transform 1 0 57224 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_622
timestamp 1666464484
transform 1 0 58328 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1666464484
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1666464484
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_27
timestamp 1666464484
transform 1 0 3588 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_31
timestamp 1666464484
transform 1 0 3956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_33
timestamp 1666464484
transform 1 0 4140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_45
timestamp 1666464484
transform 1 0 5244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_57
timestamp 1666464484
transform 1 0 6348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_69
timestamp 1666464484
transform 1 0 7452 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_81
timestamp 1666464484
transform 1 0 8556 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_93
timestamp 1666464484
transform 1 0 9660 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_98
timestamp 1666464484
transform 1 0 10120 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_110
timestamp 1666464484
transform 1 0 11224 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_122
timestamp 1666464484
transform 1 0 12328 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_134
timestamp 1666464484
transform 1 0 13432 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_146
timestamp 1666464484
transform 1 0 14536 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_158
timestamp 1666464484
transform 1 0 15640 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_163
timestamp 1666464484
transform 1 0 16100 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_175
timestamp 1666464484
transform 1 0 17204 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_187
timestamp 1666464484
transform 1 0 18308 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_199
timestamp 1666464484
transform 1 0 19412 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_211
timestamp 1666464484
transform 1 0 20516 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_223
timestamp 1666464484
transform 1 0 21620 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_228
timestamp 1666464484
transform 1 0 22080 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_240
timestamp 1666464484
transform 1 0 23184 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_252
timestamp 1666464484
transform 1 0 24288 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_264
timestamp 1666464484
transform 1 0 25392 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_276
timestamp 1666464484
transform 1 0 26496 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_288
timestamp 1666464484
transform 1 0 27600 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_293
timestamp 1666464484
transform 1 0 28060 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_305
timestamp 1666464484
transform 1 0 29164 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_317
timestamp 1666464484
transform 1 0 30268 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_329
timestamp 1666464484
transform 1 0 31372 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_341
timestamp 1666464484
transform 1 0 32476 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_353
timestamp 1666464484
transform 1 0 33580 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_358
timestamp 1666464484
transform 1 0 34040 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_370
timestamp 1666464484
transform 1 0 35144 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_382
timestamp 1666464484
transform 1 0 36248 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_394
timestamp 1666464484
transform 1 0 37352 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_406
timestamp 1666464484
transform 1 0 38456 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_418
timestamp 1666464484
transform 1 0 39560 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_423
timestamp 1666464484
transform 1 0 40020 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_435
timestamp 1666464484
transform 1 0 41124 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_447
timestamp 1666464484
transform 1 0 42228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_459
timestamp 1666464484
transform 1 0 43332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_471
timestamp 1666464484
transform 1 0 44436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_483
timestamp 1666464484
transform 1 0 45540 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_488
timestamp 1666464484
transform 1 0 46000 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_500
timestamp 1666464484
transform 1 0 47104 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_512
timestamp 1666464484
transform 1 0 48208 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_524
timestamp 1666464484
transform 1 0 49312 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_536
timestamp 1666464484
transform 1 0 50416 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_548
timestamp 1666464484
transform 1 0 51520 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_553
timestamp 1666464484
transform 1 0 51980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_565
timestamp 1666464484
transform 1 0 53084 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_577
timestamp 1666464484
transform 1 0 54188 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1666464484
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1666464484
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_613
timestamp 1666464484
transform 1 0 57500 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_618
timestamp 1666464484
transform 1 0 57960 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_624
timestamp 1666464484
transform 1 0 58512 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1666464484
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1666464484
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1666464484
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1666464484
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_51
timestamp 1666464484
transform 1 0 5796 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_63
timestamp 1666464484
transform 1 0 6900 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_66
timestamp 1666464484
transform 1 0 7176 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_78
timestamp 1666464484
transform 1 0 8280 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_90
timestamp 1666464484
transform 1 0 9384 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_102
timestamp 1666464484
transform 1 0 10488 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_114
timestamp 1666464484
transform 1 0 11592 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_126
timestamp 1666464484
transform 1 0 12696 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_131
timestamp 1666464484
transform 1 0 13156 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_143
timestamp 1666464484
transform 1 0 14260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_155
timestamp 1666464484
transform 1 0 15364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_167
timestamp 1666464484
transform 1 0 16468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_179
timestamp 1666464484
transform 1 0 17572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_191
timestamp 1666464484
transform 1 0 18676 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_196
timestamp 1666464484
transform 1 0 19136 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_208
timestamp 1666464484
transform 1 0 20240 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_220
timestamp 1666464484
transform 1 0 21344 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_232
timestamp 1666464484
transform 1 0 22448 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_244
timestamp 1666464484
transform 1 0 23552 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_256
timestamp 1666464484
transform 1 0 24656 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1666464484
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_273
timestamp 1666464484
transform 1 0 26220 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_285
timestamp 1666464484
transform 1 0 27324 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_297
timestamp 1666464484
transform 1 0 28428 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_309
timestamp 1666464484
transform 1 0 29532 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_321
timestamp 1666464484
transform 1 0 30636 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_326
timestamp 1666464484
transform 1 0 31096 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_338
timestamp 1666464484
transform 1 0 32200 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_350
timestamp 1666464484
transform 1 0 33304 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_362
timestamp 1666464484
transform 1 0 34408 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_374
timestamp 1666464484
transform 1 0 35512 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_386
timestamp 1666464484
transform 1 0 36616 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_391
timestamp 1666464484
transform 1 0 37076 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_403
timestamp 1666464484
transform 1 0 38180 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_415
timestamp 1666464484
transform 1 0 39284 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_427
timestamp 1666464484
transform 1 0 40388 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_439
timestamp 1666464484
transform 1 0 41492 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_451
timestamp 1666464484
transform 1 0 42596 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_456
timestamp 1666464484
transform 1 0 43056 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_468
timestamp 1666464484
transform 1 0 44160 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_480
timestamp 1666464484
transform 1 0 45264 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_492
timestamp 1666464484
transform 1 0 46368 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_504
timestamp 1666464484
transform 1 0 47472 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_516
timestamp 1666464484
transform 1 0 48576 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_521
timestamp 1666464484
transform 1 0 49036 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_533
timestamp 1666464484
transform 1 0 50140 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_545
timestamp 1666464484
transform 1 0 51244 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_557
timestamp 1666464484
transform 1 0 52348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_569
timestamp 1666464484
transform 1 0 53452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_581
timestamp 1666464484
transform 1 0 54556 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_586
timestamp 1666464484
transform 1 0 55016 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_598
timestamp 1666464484
transform 1 0 56120 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_610
timestamp 1666464484
transform 1 0 57224 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_622
timestamp 1666464484
transform 1 0 58328 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1666464484
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1666464484
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_27
timestamp 1666464484
transform 1 0 3588 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_31
timestamp 1666464484
transform 1 0 3956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_33
timestamp 1666464484
transform 1 0 4140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_45
timestamp 1666464484
transform 1 0 5244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_57
timestamp 1666464484
transform 1 0 6348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_69
timestamp 1666464484
transform 1 0 7452 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_81
timestamp 1666464484
transform 1 0 8556 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_93
timestamp 1666464484
transform 1 0 9660 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_98
timestamp 1666464484
transform 1 0 10120 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_110
timestamp 1666464484
transform 1 0 11224 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_122
timestamp 1666464484
transform 1 0 12328 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_134
timestamp 1666464484
transform 1 0 13432 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_146
timestamp 1666464484
transform 1 0 14536 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_158
timestamp 1666464484
transform 1 0 15640 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_163
timestamp 1666464484
transform 1 0 16100 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_175
timestamp 1666464484
transform 1 0 17204 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_187
timestamp 1666464484
transform 1 0 18308 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_199
timestamp 1666464484
transform 1 0 19412 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_211
timestamp 1666464484
transform 1 0 20516 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_223
timestamp 1666464484
transform 1 0 21620 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_228
timestamp 1666464484
transform 1 0 22080 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_240
timestamp 1666464484
transform 1 0 23184 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_252
timestamp 1666464484
transform 1 0 24288 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_264
timestamp 1666464484
transform 1 0 25392 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_276
timestamp 1666464484
transform 1 0 26496 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_288
timestamp 1666464484
transform 1 0 27600 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_293
timestamp 1666464484
transform 1 0 28060 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_305
timestamp 1666464484
transform 1 0 29164 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_317
timestamp 1666464484
transform 1 0 30268 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_329
timestamp 1666464484
transform 1 0 31372 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_341
timestamp 1666464484
transform 1 0 32476 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_353
timestamp 1666464484
transform 1 0 33580 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_358
timestamp 1666464484
transform 1 0 34040 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_370
timestamp 1666464484
transform 1 0 35144 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_382
timestamp 1666464484
transform 1 0 36248 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_394
timestamp 1666464484
transform 1 0 37352 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_406
timestamp 1666464484
transform 1 0 38456 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_418
timestamp 1666464484
transform 1 0 39560 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_423
timestamp 1666464484
transform 1 0 40020 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_435
timestamp 1666464484
transform 1 0 41124 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_447
timestamp 1666464484
transform 1 0 42228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_459
timestamp 1666464484
transform 1 0 43332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_471
timestamp 1666464484
transform 1 0 44436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_483
timestamp 1666464484
transform 1 0 45540 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_488
timestamp 1666464484
transform 1 0 46000 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_500
timestamp 1666464484
transform 1 0 47104 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_512
timestamp 1666464484
transform 1 0 48208 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_524
timestamp 1666464484
transform 1 0 49312 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_536
timestamp 1666464484
transform 1 0 50416 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_548
timestamp 1666464484
transform 1 0 51520 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_553
timestamp 1666464484
transform 1 0 51980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_565
timestamp 1666464484
transform 1 0 53084 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_577
timestamp 1666464484
transform 1 0 54188 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1666464484
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1666464484
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_613
timestamp 1666464484
transform 1 0 57500 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_618
timestamp 1666464484
transform 1 0 57960 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_624
timestamp 1666464484
transform 1 0 58512 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1666464484
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1666464484
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1666464484
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1666464484
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_51
timestamp 1666464484
transform 1 0 5796 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_63
timestamp 1666464484
transform 1 0 6900 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_66
timestamp 1666464484
transform 1 0 7176 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_78
timestamp 1666464484
transform 1 0 8280 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_90
timestamp 1666464484
transform 1 0 9384 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_102
timestamp 1666464484
transform 1 0 10488 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_114
timestamp 1666464484
transform 1 0 11592 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_126
timestamp 1666464484
transform 1 0 12696 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_131
timestamp 1666464484
transform 1 0 13156 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_143
timestamp 1666464484
transform 1 0 14260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_155
timestamp 1666464484
transform 1 0 15364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_167
timestamp 1666464484
transform 1 0 16468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_179
timestamp 1666464484
transform 1 0 17572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_191
timestamp 1666464484
transform 1 0 18676 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_196
timestamp 1666464484
transform 1 0 19136 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_208
timestamp 1666464484
transform 1 0 20240 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_220
timestamp 1666464484
transform 1 0 21344 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_232
timestamp 1666464484
transform 1 0 22448 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_244
timestamp 1666464484
transform 1 0 23552 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_256
timestamp 1666464484
transform 1 0 24656 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1666464484
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_273
timestamp 1666464484
transform 1 0 26220 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_285
timestamp 1666464484
transform 1 0 27324 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_297
timestamp 1666464484
transform 1 0 28428 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_309
timestamp 1666464484
transform 1 0 29532 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_321
timestamp 1666464484
transform 1 0 30636 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_326
timestamp 1666464484
transform 1 0 31096 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_338
timestamp 1666464484
transform 1 0 32200 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_350
timestamp 1666464484
transform 1 0 33304 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_362
timestamp 1666464484
transform 1 0 34408 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_374
timestamp 1666464484
transform 1 0 35512 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_386
timestamp 1666464484
transform 1 0 36616 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_391
timestamp 1666464484
transform 1 0 37076 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_403
timestamp 1666464484
transform 1 0 38180 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_415
timestamp 1666464484
transform 1 0 39284 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_427
timestamp 1666464484
transform 1 0 40388 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_439
timestamp 1666464484
transform 1 0 41492 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_451
timestamp 1666464484
transform 1 0 42596 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_456
timestamp 1666464484
transform 1 0 43056 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_468
timestamp 1666464484
transform 1 0 44160 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_480
timestamp 1666464484
transform 1 0 45264 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_492
timestamp 1666464484
transform 1 0 46368 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_504
timestamp 1666464484
transform 1 0 47472 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_516
timestamp 1666464484
transform 1 0 48576 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_521
timestamp 1666464484
transform 1 0 49036 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_533
timestamp 1666464484
transform 1 0 50140 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_545
timestamp 1666464484
transform 1 0 51244 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_557
timestamp 1666464484
transform 1 0 52348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_569
timestamp 1666464484
transform 1 0 53452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_581
timestamp 1666464484
transform 1 0 54556 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_586
timestamp 1666464484
transform 1 0 55016 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_598
timestamp 1666464484
transform 1 0 56120 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_610
timestamp 1666464484
transform 1 0 57224 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_622
timestamp 1666464484
transform 1 0 58328 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1666464484
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1666464484
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_27
timestamp 1666464484
transform 1 0 3588 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_31
timestamp 1666464484
transform 1 0 3956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_33
timestamp 1666464484
transform 1 0 4140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_45
timestamp 1666464484
transform 1 0 5244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_57
timestamp 1666464484
transform 1 0 6348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_69
timestamp 1666464484
transform 1 0 7452 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_81
timestamp 1666464484
transform 1 0 8556 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_93
timestamp 1666464484
transform 1 0 9660 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_98
timestamp 1666464484
transform 1 0 10120 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_110
timestamp 1666464484
transform 1 0 11224 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_122
timestamp 1666464484
transform 1 0 12328 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_134
timestamp 1666464484
transform 1 0 13432 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_146
timestamp 1666464484
transform 1 0 14536 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_158
timestamp 1666464484
transform 1 0 15640 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_163
timestamp 1666464484
transform 1 0 16100 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_175
timestamp 1666464484
transform 1 0 17204 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_187
timestamp 1666464484
transform 1 0 18308 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_199
timestamp 1666464484
transform 1 0 19412 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_211
timestamp 1666464484
transform 1 0 20516 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_223
timestamp 1666464484
transform 1 0 21620 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_228
timestamp 1666464484
transform 1 0 22080 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_240
timestamp 1666464484
transform 1 0 23184 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_252
timestamp 1666464484
transform 1 0 24288 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_264
timestamp 1666464484
transform 1 0 25392 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_276
timestamp 1666464484
transform 1 0 26496 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_288
timestamp 1666464484
transform 1 0 27600 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_293
timestamp 1666464484
transform 1 0 28060 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_305
timestamp 1666464484
transform 1 0 29164 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_317
timestamp 1666464484
transform 1 0 30268 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_329
timestamp 1666464484
transform 1 0 31372 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_341
timestamp 1666464484
transform 1 0 32476 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_353
timestamp 1666464484
transform 1 0 33580 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_358
timestamp 1666464484
transform 1 0 34040 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_370
timestamp 1666464484
transform 1 0 35144 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_382
timestamp 1666464484
transform 1 0 36248 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_394
timestamp 1666464484
transform 1 0 37352 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_406
timestamp 1666464484
transform 1 0 38456 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_418
timestamp 1666464484
transform 1 0 39560 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_423
timestamp 1666464484
transform 1 0 40020 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_435
timestamp 1666464484
transform 1 0 41124 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_447
timestamp 1666464484
transform 1 0 42228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_459
timestamp 1666464484
transform 1 0 43332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_471
timestamp 1666464484
transform 1 0 44436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_483
timestamp 1666464484
transform 1 0 45540 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_488
timestamp 1666464484
transform 1 0 46000 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_500
timestamp 1666464484
transform 1 0 47104 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_512
timestamp 1666464484
transform 1 0 48208 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_524
timestamp 1666464484
transform 1 0 49312 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_536
timestamp 1666464484
transform 1 0 50416 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_548
timestamp 1666464484
transform 1 0 51520 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_553
timestamp 1666464484
transform 1 0 51980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_565
timestamp 1666464484
transform 1 0 53084 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_577
timestamp 1666464484
transform 1 0 54188 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1666464484
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1666464484
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_613
timestamp 1666464484
transform 1 0 57500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_618
timestamp 1666464484
transform 1 0 57960 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_624
timestamp 1666464484
transform 1 0 58512 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1666464484
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1666464484
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1666464484
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1666464484
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_51
timestamp 1666464484
transform 1 0 5796 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_63
timestamp 1666464484
transform 1 0 6900 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_66
timestamp 1666464484
transform 1 0 7176 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_78
timestamp 1666464484
transform 1 0 8280 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_90
timestamp 1666464484
transform 1 0 9384 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_102
timestamp 1666464484
transform 1 0 10488 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_114
timestamp 1666464484
transform 1 0 11592 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_126
timestamp 1666464484
transform 1 0 12696 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_131
timestamp 1666464484
transform 1 0 13156 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_143
timestamp 1666464484
transform 1 0 14260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_155
timestamp 1666464484
transform 1 0 15364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_167
timestamp 1666464484
transform 1 0 16468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_179
timestamp 1666464484
transform 1 0 17572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_191
timestamp 1666464484
transform 1 0 18676 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_196
timestamp 1666464484
transform 1 0 19136 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_208
timestamp 1666464484
transform 1 0 20240 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_220
timestamp 1666464484
transform 1 0 21344 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_232
timestamp 1666464484
transform 1 0 22448 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_244
timestamp 1666464484
transform 1 0 23552 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_256
timestamp 1666464484
transform 1 0 24656 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1666464484
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_273
timestamp 1666464484
transform 1 0 26220 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_285
timestamp 1666464484
transform 1 0 27324 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_297
timestamp 1666464484
transform 1 0 28428 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_309
timestamp 1666464484
transform 1 0 29532 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_321
timestamp 1666464484
transform 1 0 30636 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_326
timestamp 1666464484
transform 1 0 31096 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_338
timestamp 1666464484
transform 1 0 32200 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_350
timestamp 1666464484
transform 1 0 33304 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_362
timestamp 1666464484
transform 1 0 34408 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_374
timestamp 1666464484
transform 1 0 35512 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_386
timestamp 1666464484
transform 1 0 36616 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_391
timestamp 1666464484
transform 1 0 37076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_403
timestamp 1666464484
transform 1 0 38180 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_415
timestamp 1666464484
transform 1 0 39284 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_427
timestamp 1666464484
transform 1 0 40388 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_439
timestamp 1666464484
transform 1 0 41492 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_451
timestamp 1666464484
transform 1 0 42596 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_456
timestamp 1666464484
transform 1 0 43056 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_468
timestamp 1666464484
transform 1 0 44160 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_480
timestamp 1666464484
transform 1 0 45264 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_492
timestamp 1666464484
transform 1 0 46368 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_504
timestamp 1666464484
transform 1 0 47472 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_516
timestamp 1666464484
transform 1 0 48576 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_521
timestamp 1666464484
transform 1 0 49036 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_533
timestamp 1666464484
transform 1 0 50140 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_545
timestamp 1666464484
transform 1 0 51244 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_557
timestamp 1666464484
transform 1 0 52348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_569
timestamp 1666464484
transform 1 0 53452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_581
timestamp 1666464484
transform 1 0 54556 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_586
timestamp 1666464484
transform 1 0 55016 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_598
timestamp 1666464484
transform 1 0 56120 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_610
timestamp 1666464484
transform 1 0 57224 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_622
timestamp 1666464484
transform 1 0 58328 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1666464484
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1666464484
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_27
timestamp 1666464484
transform 1 0 3588 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_31
timestamp 1666464484
transform 1 0 3956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_33
timestamp 1666464484
transform 1 0 4140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_45
timestamp 1666464484
transform 1 0 5244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_57
timestamp 1666464484
transform 1 0 6348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_69
timestamp 1666464484
transform 1 0 7452 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_81
timestamp 1666464484
transform 1 0 8556 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_93
timestamp 1666464484
transform 1 0 9660 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_98
timestamp 1666464484
transform 1 0 10120 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_110
timestamp 1666464484
transform 1 0 11224 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_122
timestamp 1666464484
transform 1 0 12328 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_134
timestamp 1666464484
transform 1 0 13432 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_146
timestamp 1666464484
transform 1 0 14536 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_158
timestamp 1666464484
transform 1 0 15640 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_163
timestamp 1666464484
transform 1 0 16100 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_175
timestamp 1666464484
transform 1 0 17204 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_187
timestamp 1666464484
transform 1 0 18308 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_199
timestamp 1666464484
transform 1 0 19412 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_211
timestamp 1666464484
transform 1 0 20516 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_223
timestamp 1666464484
transform 1 0 21620 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_228
timestamp 1666464484
transform 1 0 22080 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_240
timestamp 1666464484
transform 1 0 23184 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_252
timestamp 1666464484
transform 1 0 24288 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_264
timestamp 1666464484
transform 1 0 25392 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_276
timestamp 1666464484
transform 1 0 26496 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_288
timestamp 1666464484
transform 1 0 27600 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_293
timestamp 1666464484
transform 1 0 28060 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_305
timestamp 1666464484
transform 1 0 29164 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_317
timestamp 1666464484
transform 1 0 30268 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_329
timestamp 1666464484
transform 1 0 31372 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_341
timestamp 1666464484
transform 1 0 32476 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_353
timestamp 1666464484
transform 1 0 33580 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_358
timestamp 1666464484
transform 1 0 34040 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_370
timestamp 1666464484
transform 1 0 35144 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_382
timestamp 1666464484
transform 1 0 36248 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_394
timestamp 1666464484
transform 1 0 37352 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_406
timestamp 1666464484
transform 1 0 38456 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_418
timestamp 1666464484
transform 1 0 39560 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_423
timestamp 1666464484
transform 1 0 40020 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_435
timestamp 1666464484
transform 1 0 41124 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_447
timestamp 1666464484
transform 1 0 42228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_459
timestamp 1666464484
transform 1 0 43332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_471
timestamp 1666464484
transform 1 0 44436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_483
timestamp 1666464484
transform 1 0 45540 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_488
timestamp 1666464484
transform 1 0 46000 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_500
timestamp 1666464484
transform 1 0 47104 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_512
timestamp 1666464484
transform 1 0 48208 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_524
timestamp 1666464484
transform 1 0 49312 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_536
timestamp 1666464484
transform 1 0 50416 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_548
timestamp 1666464484
transform 1 0 51520 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_553
timestamp 1666464484
transform 1 0 51980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_565
timestamp 1666464484
transform 1 0 53084 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_577
timestamp 1666464484
transform 1 0 54188 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1666464484
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1666464484
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_613
timestamp 1666464484
transform 1 0 57500 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_618
timestamp 1666464484
transform 1 0 57960 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_624
timestamp 1666464484
transform 1 0 58512 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1666464484
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1666464484
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1666464484
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1666464484
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_51
timestamp 1666464484
transform 1 0 5796 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_63
timestamp 1666464484
transform 1 0 6900 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_66
timestamp 1666464484
transform 1 0 7176 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_78
timestamp 1666464484
transform 1 0 8280 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_90
timestamp 1666464484
transform 1 0 9384 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_102
timestamp 1666464484
transform 1 0 10488 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_114
timestamp 1666464484
transform 1 0 11592 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_126
timestamp 1666464484
transform 1 0 12696 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_131
timestamp 1666464484
transform 1 0 13156 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_143
timestamp 1666464484
transform 1 0 14260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_155
timestamp 1666464484
transform 1 0 15364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_167
timestamp 1666464484
transform 1 0 16468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_179
timestamp 1666464484
transform 1 0 17572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_191
timestamp 1666464484
transform 1 0 18676 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_196
timestamp 1666464484
transform 1 0 19136 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_208
timestamp 1666464484
transform 1 0 20240 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_220
timestamp 1666464484
transform 1 0 21344 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_232
timestamp 1666464484
transform 1 0 22448 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_244
timestamp 1666464484
transform 1 0 23552 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_256
timestamp 1666464484
transform 1 0 24656 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1666464484
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_273
timestamp 1666464484
transform 1 0 26220 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_285
timestamp 1666464484
transform 1 0 27324 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_297
timestamp 1666464484
transform 1 0 28428 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_309
timestamp 1666464484
transform 1 0 29532 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_321
timestamp 1666464484
transform 1 0 30636 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_326
timestamp 1666464484
transform 1 0 31096 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_338
timestamp 1666464484
transform 1 0 32200 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_350
timestamp 1666464484
transform 1 0 33304 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_362
timestamp 1666464484
transform 1 0 34408 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_374
timestamp 1666464484
transform 1 0 35512 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_386
timestamp 1666464484
transform 1 0 36616 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_391
timestamp 1666464484
transform 1 0 37076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_403
timestamp 1666464484
transform 1 0 38180 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_415
timestamp 1666464484
transform 1 0 39284 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_427
timestamp 1666464484
transform 1 0 40388 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_439
timestamp 1666464484
transform 1 0 41492 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_451
timestamp 1666464484
transform 1 0 42596 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_456
timestamp 1666464484
transform 1 0 43056 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_468
timestamp 1666464484
transform 1 0 44160 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_480
timestamp 1666464484
transform 1 0 45264 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_492
timestamp 1666464484
transform 1 0 46368 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_504
timestamp 1666464484
transform 1 0 47472 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_516
timestamp 1666464484
transform 1 0 48576 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_521
timestamp 1666464484
transform 1 0 49036 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_533
timestamp 1666464484
transform 1 0 50140 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_545
timestamp 1666464484
transform 1 0 51244 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_557
timestamp 1666464484
transform 1 0 52348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_569
timestamp 1666464484
transform 1 0 53452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_581
timestamp 1666464484
transform 1 0 54556 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_586
timestamp 1666464484
transform 1 0 55016 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_598
timestamp 1666464484
transform 1 0 56120 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_610
timestamp 1666464484
transform 1 0 57224 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_622
timestamp 1666464484
transform 1 0 58328 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1666464484
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1666464484
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_27
timestamp 1666464484
transform 1 0 3588 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_31
timestamp 1666464484
transform 1 0 3956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_33
timestamp 1666464484
transform 1 0 4140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_45
timestamp 1666464484
transform 1 0 5244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_57
timestamp 1666464484
transform 1 0 6348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_69
timestamp 1666464484
transform 1 0 7452 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_81
timestamp 1666464484
transform 1 0 8556 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_93
timestamp 1666464484
transform 1 0 9660 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_98
timestamp 1666464484
transform 1 0 10120 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_110
timestamp 1666464484
transform 1 0 11224 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_122
timestamp 1666464484
transform 1 0 12328 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_134
timestamp 1666464484
transform 1 0 13432 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_146
timestamp 1666464484
transform 1 0 14536 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_158
timestamp 1666464484
transform 1 0 15640 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_163
timestamp 1666464484
transform 1 0 16100 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_175
timestamp 1666464484
transform 1 0 17204 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_187
timestamp 1666464484
transform 1 0 18308 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_199
timestamp 1666464484
transform 1 0 19412 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_211
timestamp 1666464484
transform 1 0 20516 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_223
timestamp 1666464484
transform 1 0 21620 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_228
timestamp 1666464484
transform 1 0 22080 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_240
timestamp 1666464484
transform 1 0 23184 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_252
timestamp 1666464484
transform 1 0 24288 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_264
timestamp 1666464484
transform 1 0 25392 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_276
timestamp 1666464484
transform 1 0 26496 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_288
timestamp 1666464484
transform 1 0 27600 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_293
timestamp 1666464484
transform 1 0 28060 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_305
timestamp 1666464484
transform 1 0 29164 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_317
timestamp 1666464484
transform 1 0 30268 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_329
timestamp 1666464484
transform 1 0 31372 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_341
timestamp 1666464484
transform 1 0 32476 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_353
timestamp 1666464484
transform 1 0 33580 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_358
timestamp 1666464484
transform 1 0 34040 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_370
timestamp 1666464484
transform 1 0 35144 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_382
timestamp 1666464484
transform 1 0 36248 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_394
timestamp 1666464484
transform 1 0 37352 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_406
timestamp 1666464484
transform 1 0 38456 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_418
timestamp 1666464484
transform 1 0 39560 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_423
timestamp 1666464484
transform 1 0 40020 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_435
timestamp 1666464484
transform 1 0 41124 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_447
timestamp 1666464484
transform 1 0 42228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_459
timestamp 1666464484
transform 1 0 43332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_471
timestamp 1666464484
transform 1 0 44436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_483
timestamp 1666464484
transform 1 0 45540 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_488
timestamp 1666464484
transform 1 0 46000 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_500
timestamp 1666464484
transform 1 0 47104 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_512
timestamp 1666464484
transform 1 0 48208 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_524
timestamp 1666464484
transform 1 0 49312 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_536
timestamp 1666464484
transform 1 0 50416 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_548
timestamp 1666464484
transform 1 0 51520 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_553
timestamp 1666464484
transform 1 0 51980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_565
timestamp 1666464484
transform 1 0 53084 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_577
timestamp 1666464484
transform 1 0 54188 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1666464484
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1666464484
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_613
timestamp 1666464484
transform 1 0 57500 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_618
timestamp 1666464484
transform 1 0 57960 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_624
timestamp 1666464484
transform 1 0 58512 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1666464484
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1666464484
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1666464484
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1666464484
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_51
timestamp 1666464484
transform 1 0 5796 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_63
timestamp 1666464484
transform 1 0 6900 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_66
timestamp 1666464484
transform 1 0 7176 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_78
timestamp 1666464484
transform 1 0 8280 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_90
timestamp 1666464484
transform 1 0 9384 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_102
timestamp 1666464484
transform 1 0 10488 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_114
timestamp 1666464484
transform 1 0 11592 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_126
timestamp 1666464484
transform 1 0 12696 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_131
timestamp 1666464484
transform 1 0 13156 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_143
timestamp 1666464484
transform 1 0 14260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_155
timestamp 1666464484
transform 1 0 15364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_167
timestamp 1666464484
transform 1 0 16468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_179
timestamp 1666464484
transform 1 0 17572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_191
timestamp 1666464484
transform 1 0 18676 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_196
timestamp 1666464484
transform 1 0 19136 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_208
timestamp 1666464484
transform 1 0 20240 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_220
timestamp 1666464484
transform 1 0 21344 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_232
timestamp 1666464484
transform 1 0 22448 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_244
timestamp 1666464484
transform 1 0 23552 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_256
timestamp 1666464484
transform 1 0 24656 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1666464484
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_273
timestamp 1666464484
transform 1 0 26220 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_285
timestamp 1666464484
transform 1 0 27324 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_297
timestamp 1666464484
transform 1 0 28428 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_309
timestamp 1666464484
transform 1 0 29532 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_321
timestamp 1666464484
transform 1 0 30636 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_326
timestamp 1666464484
transform 1 0 31096 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_338
timestamp 1666464484
transform 1 0 32200 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_350
timestamp 1666464484
transform 1 0 33304 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_362
timestamp 1666464484
transform 1 0 34408 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_374
timestamp 1666464484
transform 1 0 35512 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_386
timestamp 1666464484
transform 1 0 36616 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_391
timestamp 1666464484
transform 1 0 37076 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_403
timestamp 1666464484
transform 1 0 38180 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_415
timestamp 1666464484
transform 1 0 39284 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_427
timestamp 1666464484
transform 1 0 40388 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_439
timestamp 1666464484
transform 1 0 41492 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_451
timestamp 1666464484
transform 1 0 42596 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_456
timestamp 1666464484
transform 1 0 43056 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_468
timestamp 1666464484
transform 1 0 44160 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_480
timestamp 1666464484
transform 1 0 45264 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_492
timestamp 1666464484
transform 1 0 46368 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_504
timestamp 1666464484
transform 1 0 47472 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_516
timestamp 1666464484
transform 1 0 48576 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_521
timestamp 1666464484
transform 1 0 49036 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_533
timestamp 1666464484
transform 1 0 50140 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_545
timestamp 1666464484
transform 1 0 51244 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_557
timestamp 1666464484
transform 1 0 52348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_569
timestamp 1666464484
transform 1 0 53452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_581
timestamp 1666464484
transform 1 0 54556 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_586
timestamp 1666464484
transform 1 0 55016 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_598
timestamp 1666464484
transform 1 0 56120 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_610
timestamp 1666464484
transform 1 0 57224 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_622
timestamp 1666464484
transform 1 0 58328 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1666464484
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1666464484
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_27
timestamp 1666464484
transform 1 0 3588 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_31
timestamp 1666464484
transform 1 0 3956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_33
timestamp 1666464484
transform 1 0 4140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_45
timestamp 1666464484
transform 1 0 5244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_57
timestamp 1666464484
transform 1 0 6348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_69
timestamp 1666464484
transform 1 0 7452 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_81
timestamp 1666464484
transform 1 0 8556 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_93
timestamp 1666464484
transform 1 0 9660 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_98
timestamp 1666464484
transform 1 0 10120 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_110
timestamp 1666464484
transform 1 0 11224 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_122
timestamp 1666464484
transform 1 0 12328 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_134
timestamp 1666464484
transform 1 0 13432 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_146
timestamp 1666464484
transform 1 0 14536 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_158
timestamp 1666464484
transform 1 0 15640 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_163
timestamp 1666464484
transform 1 0 16100 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_175
timestamp 1666464484
transform 1 0 17204 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_187
timestamp 1666464484
transform 1 0 18308 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_199
timestamp 1666464484
transform 1 0 19412 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_211
timestamp 1666464484
transform 1 0 20516 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_223
timestamp 1666464484
transform 1 0 21620 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_228
timestamp 1666464484
transform 1 0 22080 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_240
timestamp 1666464484
transform 1 0 23184 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_252
timestamp 1666464484
transform 1 0 24288 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_264
timestamp 1666464484
transform 1 0 25392 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_276
timestamp 1666464484
transform 1 0 26496 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_288
timestamp 1666464484
transform 1 0 27600 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_293
timestamp 1666464484
transform 1 0 28060 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_305
timestamp 1666464484
transform 1 0 29164 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_317
timestamp 1666464484
transform 1 0 30268 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_329
timestamp 1666464484
transform 1 0 31372 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_341
timestamp 1666464484
transform 1 0 32476 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_353
timestamp 1666464484
transform 1 0 33580 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_358
timestamp 1666464484
transform 1 0 34040 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_370
timestamp 1666464484
transform 1 0 35144 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_382
timestamp 1666464484
transform 1 0 36248 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_394
timestamp 1666464484
transform 1 0 37352 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_406
timestamp 1666464484
transform 1 0 38456 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_418
timestamp 1666464484
transform 1 0 39560 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_423
timestamp 1666464484
transform 1 0 40020 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_435
timestamp 1666464484
transform 1 0 41124 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_447
timestamp 1666464484
transform 1 0 42228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_459
timestamp 1666464484
transform 1 0 43332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_471
timestamp 1666464484
transform 1 0 44436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_483
timestamp 1666464484
transform 1 0 45540 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_488
timestamp 1666464484
transform 1 0 46000 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_500
timestamp 1666464484
transform 1 0 47104 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_512
timestamp 1666464484
transform 1 0 48208 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_524
timestamp 1666464484
transform 1 0 49312 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_536
timestamp 1666464484
transform 1 0 50416 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_548
timestamp 1666464484
transform 1 0 51520 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_553
timestamp 1666464484
transform 1 0 51980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_565
timestamp 1666464484
transform 1 0 53084 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_577
timestamp 1666464484
transform 1 0 54188 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1666464484
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1666464484
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_613
timestamp 1666464484
transform 1 0 57500 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_618
timestamp 1666464484
transform 1 0 57960 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_624
timestamp 1666464484
transform 1 0 58512 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1666464484
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1666464484
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1666464484
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1666464484
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_51
timestamp 1666464484
transform 1 0 5796 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_63
timestamp 1666464484
transform 1 0 6900 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_66
timestamp 1666464484
transform 1 0 7176 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_78
timestamp 1666464484
transform 1 0 8280 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_90
timestamp 1666464484
transform 1 0 9384 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_102
timestamp 1666464484
transform 1 0 10488 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_114
timestamp 1666464484
transform 1 0 11592 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_126
timestamp 1666464484
transform 1 0 12696 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_131
timestamp 1666464484
transform 1 0 13156 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_143
timestamp 1666464484
transform 1 0 14260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_155
timestamp 1666464484
transform 1 0 15364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_167
timestamp 1666464484
transform 1 0 16468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_179
timestamp 1666464484
transform 1 0 17572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_191
timestamp 1666464484
transform 1 0 18676 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_196
timestamp 1666464484
transform 1 0 19136 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_208
timestamp 1666464484
transform 1 0 20240 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_220
timestamp 1666464484
transform 1 0 21344 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_232
timestamp 1666464484
transform 1 0 22448 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_244
timestamp 1666464484
transform 1 0 23552 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_256
timestamp 1666464484
transform 1 0 24656 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1666464484
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_273
timestamp 1666464484
transform 1 0 26220 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_285
timestamp 1666464484
transform 1 0 27324 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_297
timestamp 1666464484
transform 1 0 28428 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_309
timestamp 1666464484
transform 1 0 29532 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_321
timestamp 1666464484
transform 1 0 30636 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_326
timestamp 1666464484
transform 1 0 31096 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_338
timestamp 1666464484
transform 1 0 32200 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_350
timestamp 1666464484
transform 1 0 33304 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_362
timestamp 1666464484
transform 1 0 34408 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_374
timestamp 1666464484
transform 1 0 35512 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_386
timestamp 1666464484
transform 1 0 36616 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_391
timestamp 1666464484
transform 1 0 37076 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_403
timestamp 1666464484
transform 1 0 38180 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_415
timestamp 1666464484
transform 1 0 39284 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_427
timestamp 1666464484
transform 1 0 40388 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_439
timestamp 1666464484
transform 1 0 41492 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_451
timestamp 1666464484
transform 1 0 42596 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_456
timestamp 1666464484
transform 1 0 43056 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_468
timestamp 1666464484
transform 1 0 44160 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_480
timestamp 1666464484
transform 1 0 45264 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_492
timestamp 1666464484
transform 1 0 46368 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_504
timestamp 1666464484
transform 1 0 47472 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_516
timestamp 1666464484
transform 1 0 48576 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_521
timestamp 1666464484
transform 1 0 49036 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_533
timestamp 1666464484
transform 1 0 50140 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_545
timestamp 1666464484
transform 1 0 51244 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_557
timestamp 1666464484
transform 1 0 52348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_569
timestamp 1666464484
transform 1 0 53452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_581
timestamp 1666464484
transform 1 0 54556 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_586
timestamp 1666464484
transform 1 0 55016 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_598
timestamp 1666464484
transform 1 0 56120 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_610
timestamp 1666464484
transform 1 0 57224 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_622
timestamp 1666464484
transform 1 0 58328 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1666464484
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1666464484
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_27
timestamp 1666464484
transform 1 0 3588 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_31
timestamp 1666464484
transform 1 0 3956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_33
timestamp 1666464484
transform 1 0 4140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_45
timestamp 1666464484
transform 1 0 5244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_57
timestamp 1666464484
transform 1 0 6348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_69
timestamp 1666464484
transform 1 0 7452 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_81
timestamp 1666464484
transform 1 0 8556 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_93
timestamp 1666464484
transform 1 0 9660 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_98
timestamp 1666464484
transform 1 0 10120 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_110
timestamp 1666464484
transform 1 0 11224 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_122
timestamp 1666464484
transform 1 0 12328 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_134
timestamp 1666464484
transform 1 0 13432 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_146
timestamp 1666464484
transform 1 0 14536 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_158
timestamp 1666464484
transform 1 0 15640 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_163
timestamp 1666464484
transform 1 0 16100 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_175
timestamp 1666464484
transform 1 0 17204 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_187
timestamp 1666464484
transform 1 0 18308 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_199
timestamp 1666464484
transform 1 0 19412 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_211
timestamp 1666464484
transform 1 0 20516 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_223
timestamp 1666464484
transform 1 0 21620 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_228
timestamp 1666464484
transform 1 0 22080 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_240
timestamp 1666464484
transform 1 0 23184 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_252
timestamp 1666464484
transform 1 0 24288 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_264
timestamp 1666464484
transform 1 0 25392 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_276
timestamp 1666464484
transform 1 0 26496 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_288
timestamp 1666464484
transform 1 0 27600 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_293
timestamp 1666464484
transform 1 0 28060 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_305
timestamp 1666464484
transform 1 0 29164 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_317
timestamp 1666464484
transform 1 0 30268 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_329
timestamp 1666464484
transform 1 0 31372 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_341
timestamp 1666464484
transform 1 0 32476 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_353
timestamp 1666464484
transform 1 0 33580 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_358
timestamp 1666464484
transform 1 0 34040 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_370
timestamp 1666464484
transform 1 0 35144 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_382
timestamp 1666464484
transform 1 0 36248 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_394
timestamp 1666464484
transform 1 0 37352 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_406
timestamp 1666464484
transform 1 0 38456 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_418
timestamp 1666464484
transform 1 0 39560 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_423
timestamp 1666464484
transform 1 0 40020 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_435
timestamp 1666464484
transform 1 0 41124 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_447
timestamp 1666464484
transform 1 0 42228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_459
timestamp 1666464484
transform 1 0 43332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_471
timestamp 1666464484
transform 1 0 44436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_483
timestamp 1666464484
transform 1 0 45540 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_488
timestamp 1666464484
transform 1 0 46000 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_500
timestamp 1666464484
transform 1 0 47104 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_512
timestamp 1666464484
transform 1 0 48208 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_524
timestamp 1666464484
transform 1 0 49312 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_536
timestamp 1666464484
transform 1 0 50416 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_548
timestamp 1666464484
transform 1 0 51520 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_553
timestamp 1666464484
transform 1 0 51980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_565
timestamp 1666464484
transform 1 0 53084 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_577
timestamp 1666464484
transform 1 0 54188 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1666464484
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1666464484
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_613
timestamp 1666464484
transform 1 0 57500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_618
timestamp 1666464484
transform 1 0 57960 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_624
timestamp 1666464484
transform 1 0 58512 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1666464484
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1666464484
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1666464484
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1666464484
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_51
timestamp 1666464484
transform 1 0 5796 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_63
timestamp 1666464484
transform 1 0 6900 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_66
timestamp 1666464484
transform 1 0 7176 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_78
timestamp 1666464484
transform 1 0 8280 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_90
timestamp 1666464484
transform 1 0 9384 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_102
timestamp 1666464484
transform 1 0 10488 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_114
timestamp 1666464484
transform 1 0 11592 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_126
timestamp 1666464484
transform 1 0 12696 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_131
timestamp 1666464484
transform 1 0 13156 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_143
timestamp 1666464484
transform 1 0 14260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_155
timestamp 1666464484
transform 1 0 15364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_167
timestamp 1666464484
transform 1 0 16468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_179
timestamp 1666464484
transform 1 0 17572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_191
timestamp 1666464484
transform 1 0 18676 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_196
timestamp 1666464484
transform 1 0 19136 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_208
timestamp 1666464484
transform 1 0 20240 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_220
timestamp 1666464484
transform 1 0 21344 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_232
timestamp 1666464484
transform 1 0 22448 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_244
timestamp 1666464484
transform 1 0 23552 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_256
timestamp 1666464484
transform 1 0 24656 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1666464484
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_273
timestamp 1666464484
transform 1 0 26220 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_285
timestamp 1666464484
transform 1 0 27324 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_297
timestamp 1666464484
transform 1 0 28428 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_309
timestamp 1666464484
transform 1 0 29532 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_321
timestamp 1666464484
transform 1 0 30636 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_326
timestamp 1666464484
transform 1 0 31096 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_338
timestamp 1666464484
transform 1 0 32200 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_350
timestamp 1666464484
transform 1 0 33304 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_362
timestamp 1666464484
transform 1 0 34408 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_374
timestamp 1666464484
transform 1 0 35512 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_386
timestamp 1666464484
transform 1 0 36616 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_391
timestamp 1666464484
transform 1 0 37076 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_403
timestamp 1666464484
transform 1 0 38180 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_415
timestamp 1666464484
transform 1 0 39284 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_427
timestamp 1666464484
transform 1 0 40388 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_439
timestamp 1666464484
transform 1 0 41492 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_451
timestamp 1666464484
transform 1 0 42596 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_456
timestamp 1666464484
transform 1 0 43056 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_468
timestamp 1666464484
transform 1 0 44160 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_480
timestamp 1666464484
transform 1 0 45264 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_492
timestamp 1666464484
transform 1 0 46368 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_504
timestamp 1666464484
transform 1 0 47472 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_516
timestamp 1666464484
transform 1 0 48576 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_521
timestamp 1666464484
transform 1 0 49036 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_533
timestamp 1666464484
transform 1 0 50140 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_545
timestamp 1666464484
transform 1 0 51244 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_557
timestamp 1666464484
transform 1 0 52348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_569
timestamp 1666464484
transform 1 0 53452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_581
timestamp 1666464484
transform 1 0 54556 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_586
timestamp 1666464484
transform 1 0 55016 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_598
timestamp 1666464484
transform 1 0 56120 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_610
timestamp 1666464484
transform 1 0 57224 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_622
timestamp 1666464484
transform 1 0 58328 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1666464484
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1666464484
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_27
timestamp 1666464484
transform 1 0 3588 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_31
timestamp 1666464484
transform 1 0 3956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_33
timestamp 1666464484
transform 1 0 4140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_45
timestamp 1666464484
transform 1 0 5244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_57
timestamp 1666464484
transform 1 0 6348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_69
timestamp 1666464484
transform 1 0 7452 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_81
timestamp 1666464484
transform 1 0 8556 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_93
timestamp 1666464484
transform 1 0 9660 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_98
timestamp 1666464484
transform 1 0 10120 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_110
timestamp 1666464484
transform 1 0 11224 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_122
timestamp 1666464484
transform 1 0 12328 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_134
timestamp 1666464484
transform 1 0 13432 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_146
timestamp 1666464484
transform 1 0 14536 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_158
timestamp 1666464484
transform 1 0 15640 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_163
timestamp 1666464484
transform 1 0 16100 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_175
timestamp 1666464484
transform 1 0 17204 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_187
timestamp 1666464484
transform 1 0 18308 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_199
timestamp 1666464484
transform 1 0 19412 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_211
timestamp 1666464484
transform 1 0 20516 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_223
timestamp 1666464484
transform 1 0 21620 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_228
timestamp 1666464484
transform 1 0 22080 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_240
timestamp 1666464484
transform 1 0 23184 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_252
timestamp 1666464484
transform 1 0 24288 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_264
timestamp 1666464484
transform 1 0 25392 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_276
timestamp 1666464484
transform 1 0 26496 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_288
timestamp 1666464484
transform 1 0 27600 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_293
timestamp 1666464484
transform 1 0 28060 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_305
timestamp 1666464484
transform 1 0 29164 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_317
timestamp 1666464484
transform 1 0 30268 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_329
timestamp 1666464484
transform 1 0 31372 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_341
timestamp 1666464484
transform 1 0 32476 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_353
timestamp 1666464484
transform 1 0 33580 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_358
timestamp 1666464484
transform 1 0 34040 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_370
timestamp 1666464484
transform 1 0 35144 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_382
timestamp 1666464484
transform 1 0 36248 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_394
timestamp 1666464484
transform 1 0 37352 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_406
timestamp 1666464484
transform 1 0 38456 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_418
timestamp 1666464484
transform 1 0 39560 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_423
timestamp 1666464484
transform 1 0 40020 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_435
timestamp 1666464484
transform 1 0 41124 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_447
timestamp 1666464484
transform 1 0 42228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_459
timestamp 1666464484
transform 1 0 43332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_471
timestamp 1666464484
transform 1 0 44436 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_483
timestamp 1666464484
transform 1 0 45540 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_488
timestamp 1666464484
transform 1 0 46000 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_500
timestamp 1666464484
transform 1 0 47104 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_512
timestamp 1666464484
transform 1 0 48208 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_524
timestamp 1666464484
transform 1 0 49312 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_536
timestamp 1666464484
transform 1 0 50416 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_548
timestamp 1666464484
transform 1 0 51520 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_553
timestamp 1666464484
transform 1 0 51980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_565
timestamp 1666464484
transform 1 0 53084 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_577
timestamp 1666464484
transform 1 0 54188 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1666464484
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1666464484
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_613
timestamp 1666464484
transform 1 0 57500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_618
timestamp 1666464484
transform 1 0 57960 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_624
timestamp 1666464484
transform 1 0 58512 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1666464484
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1666464484
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1666464484
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1666464484
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_51
timestamp 1666464484
transform 1 0 5796 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_63
timestamp 1666464484
transform 1 0 6900 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_66
timestamp 1666464484
transform 1 0 7176 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_78
timestamp 1666464484
transform 1 0 8280 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_90
timestamp 1666464484
transform 1 0 9384 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_102
timestamp 1666464484
transform 1 0 10488 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_114
timestamp 1666464484
transform 1 0 11592 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_126
timestamp 1666464484
transform 1 0 12696 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_131
timestamp 1666464484
transform 1 0 13156 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_143
timestamp 1666464484
transform 1 0 14260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_155
timestamp 1666464484
transform 1 0 15364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_167
timestamp 1666464484
transform 1 0 16468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_179
timestamp 1666464484
transform 1 0 17572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_191
timestamp 1666464484
transform 1 0 18676 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_196
timestamp 1666464484
transform 1 0 19136 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_208
timestamp 1666464484
transform 1 0 20240 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_220
timestamp 1666464484
transform 1 0 21344 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_232
timestamp 1666464484
transform 1 0 22448 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_244
timestamp 1666464484
transform 1 0 23552 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_256
timestamp 1666464484
transform 1 0 24656 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1666464484
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_273
timestamp 1666464484
transform 1 0 26220 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_285
timestamp 1666464484
transform 1 0 27324 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_297
timestamp 1666464484
transform 1 0 28428 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_309
timestamp 1666464484
transform 1 0 29532 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_321
timestamp 1666464484
transform 1 0 30636 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_326
timestamp 1666464484
transform 1 0 31096 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_338
timestamp 1666464484
transform 1 0 32200 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_350
timestamp 1666464484
transform 1 0 33304 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_362
timestamp 1666464484
transform 1 0 34408 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_374
timestamp 1666464484
transform 1 0 35512 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_386
timestamp 1666464484
transform 1 0 36616 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_391
timestamp 1666464484
transform 1 0 37076 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_403
timestamp 1666464484
transform 1 0 38180 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_415
timestamp 1666464484
transform 1 0 39284 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_427
timestamp 1666464484
transform 1 0 40388 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_439
timestamp 1666464484
transform 1 0 41492 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_451
timestamp 1666464484
transform 1 0 42596 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_456
timestamp 1666464484
transform 1 0 43056 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_468
timestamp 1666464484
transform 1 0 44160 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_480
timestamp 1666464484
transform 1 0 45264 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_492
timestamp 1666464484
transform 1 0 46368 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_504
timestamp 1666464484
transform 1 0 47472 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_516
timestamp 1666464484
transform 1 0 48576 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_521
timestamp 1666464484
transform 1 0 49036 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_533
timestamp 1666464484
transform 1 0 50140 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_545
timestamp 1666464484
transform 1 0 51244 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_557
timestamp 1666464484
transform 1 0 52348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_569
timestamp 1666464484
transform 1 0 53452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_581
timestamp 1666464484
transform 1 0 54556 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_586
timestamp 1666464484
transform 1 0 55016 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_598
timestamp 1666464484
transform 1 0 56120 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_610
timestamp 1666464484
transform 1 0 57224 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_622
timestamp 1666464484
transform 1 0 58328 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1666464484
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1666464484
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_27
timestamp 1666464484
transform 1 0 3588 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_31
timestamp 1666464484
transform 1 0 3956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_33
timestamp 1666464484
transform 1 0 4140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_45
timestamp 1666464484
transform 1 0 5244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_57
timestamp 1666464484
transform 1 0 6348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_69
timestamp 1666464484
transform 1 0 7452 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_81
timestamp 1666464484
transform 1 0 8556 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_93
timestamp 1666464484
transform 1 0 9660 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_98
timestamp 1666464484
transform 1 0 10120 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_110
timestamp 1666464484
transform 1 0 11224 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_122
timestamp 1666464484
transform 1 0 12328 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_134
timestamp 1666464484
transform 1 0 13432 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_146
timestamp 1666464484
transform 1 0 14536 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_158
timestamp 1666464484
transform 1 0 15640 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_163
timestamp 1666464484
transform 1 0 16100 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_175
timestamp 1666464484
transform 1 0 17204 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_187
timestamp 1666464484
transform 1 0 18308 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_199
timestamp 1666464484
transform 1 0 19412 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_211
timestamp 1666464484
transform 1 0 20516 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_223
timestamp 1666464484
transform 1 0 21620 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_228
timestamp 1666464484
transform 1 0 22080 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_240
timestamp 1666464484
transform 1 0 23184 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_252
timestamp 1666464484
transform 1 0 24288 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_264
timestamp 1666464484
transform 1 0 25392 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_276
timestamp 1666464484
transform 1 0 26496 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_288
timestamp 1666464484
transform 1 0 27600 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_293
timestamp 1666464484
transform 1 0 28060 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_305
timestamp 1666464484
transform 1 0 29164 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_317
timestamp 1666464484
transform 1 0 30268 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_329
timestamp 1666464484
transform 1 0 31372 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_341
timestamp 1666464484
transform 1 0 32476 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_353
timestamp 1666464484
transform 1 0 33580 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_358
timestamp 1666464484
transform 1 0 34040 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_370
timestamp 1666464484
transform 1 0 35144 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_382
timestamp 1666464484
transform 1 0 36248 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_394
timestamp 1666464484
transform 1 0 37352 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_406
timestamp 1666464484
transform 1 0 38456 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_418
timestamp 1666464484
transform 1 0 39560 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_423
timestamp 1666464484
transform 1 0 40020 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_435
timestamp 1666464484
transform 1 0 41124 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_447
timestamp 1666464484
transform 1 0 42228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_459
timestamp 1666464484
transform 1 0 43332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_471
timestamp 1666464484
transform 1 0 44436 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_483
timestamp 1666464484
transform 1 0 45540 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_488
timestamp 1666464484
transform 1 0 46000 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_500
timestamp 1666464484
transform 1 0 47104 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_512
timestamp 1666464484
transform 1 0 48208 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_524
timestamp 1666464484
transform 1 0 49312 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_536
timestamp 1666464484
transform 1 0 50416 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_548
timestamp 1666464484
transform 1 0 51520 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_553
timestamp 1666464484
transform 1 0 51980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_565
timestamp 1666464484
transform 1 0 53084 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_577
timestamp 1666464484
transform 1 0 54188 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1666464484
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1666464484
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_613
timestamp 1666464484
transform 1 0 57500 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_618
timestamp 1666464484
transform 1 0 57960 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_624
timestamp 1666464484
transform 1 0 58512 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1666464484
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1666464484
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1666464484
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1666464484
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_51
timestamp 1666464484
transform 1 0 5796 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_63
timestamp 1666464484
transform 1 0 6900 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_66
timestamp 1666464484
transform 1 0 7176 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_78
timestamp 1666464484
transform 1 0 8280 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_90
timestamp 1666464484
transform 1 0 9384 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_102
timestamp 1666464484
transform 1 0 10488 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_114
timestamp 1666464484
transform 1 0 11592 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_126
timestamp 1666464484
transform 1 0 12696 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_131
timestamp 1666464484
transform 1 0 13156 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_143
timestamp 1666464484
transform 1 0 14260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_155
timestamp 1666464484
transform 1 0 15364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_167
timestamp 1666464484
transform 1 0 16468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_179
timestamp 1666464484
transform 1 0 17572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_191
timestamp 1666464484
transform 1 0 18676 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_196
timestamp 1666464484
transform 1 0 19136 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_208
timestamp 1666464484
transform 1 0 20240 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_220
timestamp 1666464484
transform 1 0 21344 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_232
timestamp 1666464484
transform 1 0 22448 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_244
timestamp 1666464484
transform 1 0 23552 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_256
timestamp 1666464484
transform 1 0 24656 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1666464484
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_273
timestamp 1666464484
transform 1 0 26220 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_285
timestamp 1666464484
transform 1 0 27324 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_297
timestamp 1666464484
transform 1 0 28428 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_309
timestamp 1666464484
transform 1 0 29532 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_321
timestamp 1666464484
transform 1 0 30636 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_326
timestamp 1666464484
transform 1 0 31096 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_338
timestamp 1666464484
transform 1 0 32200 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_350
timestamp 1666464484
transform 1 0 33304 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_362
timestamp 1666464484
transform 1 0 34408 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_374
timestamp 1666464484
transform 1 0 35512 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_386
timestamp 1666464484
transform 1 0 36616 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_391
timestamp 1666464484
transform 1 0 37076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_403
timestamp 1666464484
transform 1 0 38180 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_415
timestamp 1666464484
transform 1 0 39284 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_427
timestamp 1666464484
transform 1 0 40388 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_439
timestamp 1666464484
transform 1 0 41492 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_451
timestamp 1666464484
transform 1 0 42596 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_456
timestamp 1666464484
transform 1 0 43056 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_468
timestamp 1666464484
transform 1 0 44160 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_480
timestamp 1666464484
transform 1 0 45264 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_492
timestamp 1666464484
transform 1 0 46368 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_504
timestamp 1666464484
transform 1 0 47472 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_516
timestamp 1666464484
transform 1 0 48576 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_521
timestamp 1666464484
transform 1 0 49036 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_533
timestamp 1666464484
transform 1 0 50140 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_545
timestamp 1666464484
transform 1 0 51244 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_557
timestamp 1666464484
transform 1 0 52348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_569
timestamp 1666464484
transform 1 0 53452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_581
timestamp 1666464484
transform 1 0 54556 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_586
timestamp 1666464484
transform 1 0 55016 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_598
timestamp 1666464484
transform 1 0 56120 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_610
timestamp 1666464484
transform 1 0 57224 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_622
timestamp 1666464484
transform 1 0 58328 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1666464484
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1666464484
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_27
timestamp 1666464484
transform 1 0 3588 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_31
timestamp 1666464484
transform 1 0 3956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_33
timestamp 1666464484
transform 1 0 4140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_45
timestamp 1666464484
transform 1 0 5244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_57
timestamp 1666464484
transform 1 0 6348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_69
timestamp 1666464484
transform 1 0 7452 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_81
timestamp 1666464484
transform 1 0 8556 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_93
timestamp 1666464484
transform 1 0 9660 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_98
timestamp 1666464484
transform 1 0 10120 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_110
timestamp 1666464484
transform 1 0 11224 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_122
timestamp 1666464484
transform 1 0 12328 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_134
timestamp 1666464484
transform 1 0 13432 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_146
timestamp 1666464484
transform 1 0 14536 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_158
timestamp 1666464484
transform 1 0 15640 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_163
timestamp 1666464484
transform 1 0 16100 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_175
timestamp 1666464484
transform 1 0 17204 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_187
timestamp 1666464484
transform 1 0 18308 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_199
timestamp 1666464484
transform 1 0 19412 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_211
timestamp 1666464484
transform 1 0 20516 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_223
timestamp 1666464484
transform 1 0 21620 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_228
timestamp 1666464484
transform 1 0 22080 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_240
timestamp 1666464484
transform 1 0 23184 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_252
timestamp 1666464484
transform 1 0 24288 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_264
timestamp 1666464484
transform 1 0 25392 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_276
timestamp 1666464484
transform 1 0 26496 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_288
timestamp 1666464484
transform 1 0 27600 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_293
timestamp 1666464484
transform 1 0 28060 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_305
timestamp 1666464484
transform 1 0 29164 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_317
timestamp 1666464484
transform 1 0 30268 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_329
timestamp 1666464484
transform 1 0 31372 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_341
timestamp 1666464484
transform 1 0 32476 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_353
timestamp 1666464484
transform 1 0 33580 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_358
timestamp 1666464484
transform 1 0 34040 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_370
timestamp 1666464484
transform 1 0 35144 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_382
timestamp 1666464484
transform 1 0 36248 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_394
timestamp 1666464484
transform 1 0 37352 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_406
timestamp 1666464484
transform 1 0 38456 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_418
timestamp 1666464484
transform 1 0 39560 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_423
timestamp 1666464484
transform 1 0 40020 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_435
timestamp 1666464484
transform 1 0 41124 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_447
timestamp 1666464484
transform 1 0 42228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_459
timestamp 1666464484
transform 1 0 43332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_471
timestamp 1666464484
transform 1 0 44436 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_483
timestamp 1666464484
transform 1 0 45540 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_488
timestamp 1666464484
transform 1 0 46000 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_500
timestamp 1666464484
transform 1 0 47104 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_512
timestamp 1666464484
transform 1 0 48208 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_524
timestamp 1666464484
transform 1 0 49312 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_536
timestamp 1666464484
transform 1 0 50416 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_548
timestamp 1666464484
transform 1 0 51520 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_553
timestamp 1666464484
transform 1 0 51980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_565
timestamp 1666464484
transform 1 0 53084 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_577
timestamp 1666464484
transform 1 0 54188 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1666464484
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1666464484
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_613
timestamp 1666464484
transform 1 0 57500 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_618
timestamp 1666464484
transform 1 0 57960 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_624
timestamp 1666464484
transform 1 0 58512 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1666464484
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1666464484
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1666464484
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1666464484
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_51
timestamp 1666464484
transform 1 0 5796 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_63
timestamp 1666464484
transform 1 0 6900 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_66
timestamp 1666464484
transform 1 0 7176 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_78
timestamp 1666464484
transform 1 0 8280 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_90
timestamp 1666464484
transform 1 0 9384 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_102
timestamp 1666464484
transform 1 0 10488 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_114
timestamp 1666464484
transform 1 0 11592 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_126
timestamp 1666464484
transform 1 0 12696 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_131
timestamp 1666464484
transform 1 0 13156 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_143
timestamp 1666464484
transform 1 0 14260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_155
timestamp 1666464484
transform 1 0 15364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_167
timestamp 1666464484
transform 1 0 16468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_179
timestamp 1666464484
transform 1 0 17572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_191
timestamp 1666464484
transform 1 0 18676 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_196
timestamp 1666464484
transform 1 0 19136 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_208
timestamp 1666464484
transform 1 0 20240 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_220
timestamp 1666464484
transform 1 0 21344 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_232
timestamp 1666464484
transform 1 0 22448 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_244
timestamp 1666464484
transform 1 0 23552 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_256
timestamp 1666464484
transform 1 0 24656 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1666464484
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_273
timestamp 1666464484
transform 1 0 26220 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_285
timestamp 1666464484
transform 1 0 27324 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_297
timestamp 1666464484
transform 1 0 28428 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_309
timestamp 1666464484
transform 1 0 29532 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_321
timestamp 1666464484
transform 1 0 30636 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_326
timestamp 1666464484
transform 1 0 31096 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_338
timestamp 1666464484
transform 1 0 32200 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_350
timestamp 1666464484
transform 1 0 33304 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_362
timestamp 1666464484
transform 1 0 34408 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_374
timestamp 1666464484
transform 1 0 35512 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_386
timestamp 1666464484
transform 1 0 36616 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_391
timestamp 1666464484
transform 1 0 37076 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_403
timestamp 1666464484
transform 1 0 38180 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_415
timestamp 1666464484
transform 1 0 39284 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_427
timestamp 1666464484
transform 1 0 40388 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_439
timestamp 1666464484
transform 1 0 41492 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_451
timestamp 1666464484
transform 1 0 42596 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_456
timestamp 1666464484
transform 1 0 43056 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_468
timestamp 1666464484
transform 1 0 44160 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_480
timestamp 1666464484
transform 1 0 45264 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_492
timestamp 1666464484
transform 1 0 46368 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_504
timestamp 1666464484
transform 1 0 47472 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_516
timestamp 1666464484
transform 1 0 48576 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_521
timestamp 1666464484
transform 1 0 49036 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_533
timestamp 1666464484
transform 1 0 50140 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_545
timestamp 1666464484
transform 1 0 51244 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_557
timestamp 1666464484
transform 1 0 52348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_569
timestamp 1666464484
transform 1 0 53452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_581
timestamp 1666464484
transform 1 0 54556 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_586
timestamp 1666464484
transform 1 0 55016 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_598
timestamp 1666464484
transform 1 0 56120 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_610
timestamp 1666464484
transform 1 0 57224 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_622
timestamp 1666464484
transform 1 0 58328 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1666464484
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1666464484
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_27
timestamp 1666464484
transform 1 0 3588 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_31
timestamp 1666464484
transform 1 0 3956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_33
timestamp 1666464484
transform 1 0 4140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_45
timestamp 1666464484
transform 1 0 5244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_57
timestamp 1666464484
transform 1 0 6348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_69
timestamp 1666464484
transform 1 0 7452 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_81
timestamp 1666464484
transform 1 0 8556 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_93
timestamp 1666464484
transform 1 0 9660 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_98
timestamp 1666464484
transform 1 0 10120 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_110
timestamp 1666464484
transform 1 0 11224 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_122
timestamp 1666464484
transform 1 0 12328 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_134
timestamp 1666464484
transform 1 0 13432 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_146
timestamp 1666464484
transform 1 0 14536 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_158
timestamp 1666464484
transform 1 0 15640 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_163
timestamp 1666464484
transform 1 0 16100 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_175
timestamp 1666464484
transform 1 0 17204 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_187
timestamp 1666464484
transform 1 0 18308 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_199
timestamp 1666464484
transform 1 0 19412 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_211
timestamp 1666464484
transform 1 0 20516 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_223
timestamp 1666464484
transform 1 0 21620 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_228
timestamp 1666464484
transform 1 0 22080 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_240
timestamp 1666464484
transform 1 0 23184 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_252
timestamp 1666464484
transform 1 0 24288 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_264
timestamp 1666464484
transform 1 0 25392 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_276
timestamp 1666464484
transform 1 0 26496 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_288
timestamp 1666464484
transform 1 0 27600 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_293
timestamp 1666464484
transform 1 0 28060 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_305
timestamp 1666464484
transform 1 0 29164 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_317
timestamp 1666464484
transform 1 0 30268 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_329
timestamp 1666464484
transform 1 0 31372 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_341
timestamp 1666464484
transform 1 0 32476 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_353
timestamp 1666464484
transform 1 0 33580 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_358
timestamp 1666464484
transform 1 0 34040 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_370
timestamp 1666464484
transform 1 0 35144 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_382
timestamp 1666464484
transform 1 0 36248 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_394
timestamp 1666464484
transform 1 0 37352 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_406
timestamp 1666464484
transform 1 0 38456 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_418
timestamp 1666464484
transform 1 0 39560 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_423
timestamp 1666464484
transform 1 0 40020 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_435
timestamp 1666464484
transform 1 0 41124 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_447
timestamp 1666464484
transform 1 0 42228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_459
timestamp 1666464484
transform 1 0 43332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_471
timestamp 1666464484
transform 1 0 44436 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_483
timestamp 1666464484
transform 1 0 45540 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_488
timestamp 1666464484
transform 1 0 46000 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_500
timestamp 1666464484
transform 1 0 47104 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_512
timestamp 1666464484
transform 1 0 48208 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_524
timestamp 1666464484
transform 1 0 49312 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_536
timestamp 1666464484
transform 1 0 50416 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_548
timestamp 1666464484
transform 1 0 51520 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_553
timestamp 1666464484
transform 1 0 51980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_565
timestamp 1666464484
transform 1 0 53084 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_577
timestamp 1666464484
transform 1 0 54188 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1666464484
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1666464484
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_613
timestamp 1666464484
transform 1 0 57500 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_88_618
timestamp 1666464484
transform 1 0 57960 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_624
timestamp 1666464484
transform 1 0 58512 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1666464484
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1666464484
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1666464484
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1666464484
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_51
timestamp 1666464484
transform 1 0 5796 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_63
timestamp 1666464484
transform 1 0 6900 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_66
timestamp 1666464484
transform 1 0 7176 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_78
timestamp 1666464484
transform 1 0 8280 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_90
timestamp 1666464484
transform 1 0 9384 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_102
timestamp 1666464484
transform 1 0 10488 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_114
timestamp 1666464484
transform 1 0 11592 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_126
timestamp 1666464484
transform 1 0 12696 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_131
timestamp 1666464484
transform 1 0 13156 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_143
timestamp 1666464484
transform 1 0 14260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_155
timestamp 1666464484
transform 1 0 15364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_167
timestamp 1666464484
transform 1 0 16468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_179
timestamp 1666464484
transform 1 0 17572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_191
timestamp 1666464484
transform 1 0 18676 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_196
timestamp 1666464484
transform 1 0 19136 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_208
timestamp 1666464484
transform 1 0 20240 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_220
timestamp 1666464484
transform 1 0 21344 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_232
timestamp 1666464484
transform 1 0 22448 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_244
timestamp 1666464484
transform 1 0 23552 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_256
timestamp 1666464484
transform 1 0 24656 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1666464484
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_273
timestamp 1666464484
transform 1 0 26220 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_285
timestamp 1666464484
transform 1 0 27324 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_297
timestamp 1666464484
transform 1 0 28428 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_309
timestamp 1666464484
transform 1 0 29532 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_321
timestamp 1666464484
transform 1 0 30636 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_326
timestamp 1666464484
transform 1 0 31096 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_338
timestamp 1666464484
transform 1 0 32200 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_350
timestamp 1666464484
transform 1 0 33304 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_362
timestamp 1666464484
transform 1 0 34408 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_374
timestamp 1666464484
transform 1 0 35512 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_386
timestamp 1666464484
transform 1 0 36616 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_391
timestamp 1666464484
transform 1 0 37076 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_403
timestamp 1666464484
transform 1 0 38180 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_415
timestamp 1666464484
transform 1 0 39284 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_427
timestamp 1666464484
transform 1 0 40388 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_439
timestamp 1666464484
transform 1 0 41492 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_451
timestamp 1666464484
transform 1 0 42596 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_456
timestamp 1666464484
transform 1 0 43056 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_468
timestamp 1666464484
transform 1 0 44160 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_480
timestamp 1666464484
transform 1 0 45264 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_492
timestamp 1666464484
transform 1 0 46368 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_504
timestamp 1666464484
transform 1 0 47472 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_516
timestamp 1666464484
transform 1 0 48576 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_521
timestamp 1666464484
transform 1 0 49036 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_533
timestamp 1666464484
transform 1 0 50140 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_545
timestamp 1666464484
transform 1 0 51244 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_557
timestamp 1666464484
transform 1 0 52348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_569
timestamp 1666464484
transform 1 0 53452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_581
timestamp 1666464484
transform 1 0 54556 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_586
timestamp 1666464484
transform 1 0 55016 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_598
timestamp 1666464484
transform 1 0 56120 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_610
timestamp 1666464484
transform 1 0 57224 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_622
timestamp 1666464484
transform 1 0 58328 0 -1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1666464484
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1666464484
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_27
timestamp 1666464484
transform 1 0 3588 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_31
timestamp 1666464484
transform 1 0 3956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_33
timestamp 1666464484
transform 1 0 4140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_45
timestamp 1666464484
transform 1 0 5244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_57
timestamp 1666464484
transform 1 0 6348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_69
timestamp 1666464484
transform 1 0 7452 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_81
timestamp 1666464484
transform 1 0 8556 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_93
timestamp 1666464484
transform 1 0 9660 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_98
timestamp 1666464484
transform 1 0 10120 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_110
timestamp 1666464484
transform 1 0 11224 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_122
timestamp 1666464484
transform 1 0 12328 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_134
timestamp 1666464484
transform 1 0 13432 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_146
timestamp 1666464484
transform 1 0 14536 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_158
timestamp 1666464484
transform 1 0 15640 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_163
timestamp 1666464484
transform 1 0 16100 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_175
timestamp 1666464484
transform 1 0 17204 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_187
timestamp 1666464484
transform 1 0 18308 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_199
timestamp 1666464484
transform 1 0 19412 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_211
timestamp 1666464484
transform 1 0 20516 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_223
timestamp 1666464484
transform 1 0 21620 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_228
timestamp 1666464484
transform 1 0 22080 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_240
timestamp 1666464484
transform 1 0 23184 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_252
timestamp 1666464484
transform 1 0 24288 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_264
timestamp 1666464484
transform 1 0 25392 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_276
timestamp 1666464484
transform 1 0 26496 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_288
timestamp 1666464484
transform 1 0 27600 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_293
timestamp 1666464484
transform 1 0 28060 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_305
timestamp 1666464484
transform 1 0 29164 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_317
timestamp 1666464484
transform 1 0 30268 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_329
timestamp 1666464484
transform 1 0 31372 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_341
timestamp 1666464484
transform 1 0 32476 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_353
timestamp 1666464484
transform 1 0 33580 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_358
timestamp 1666464484
transform 1 0 34040 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_363
timestamp 1666464484
transform 1 0 34500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_375
timestamp 1666464484
transform 1 0 35604 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_387
timestamp 1666464484
transform 1 0 36708 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_399
timestamp 1666464484
transform 1 0 37812 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_411
timestamp 1666464484
transform 1 0 38916 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_90_419
timestamp 1666464484
transform 1 0 39652 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_423
timestamp 1666464484
transform 1 0 40020 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_435
timestamp 1666464484
transform 1 0 41124 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_447
timestamp 1666464484
transform 1 0 42228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_459
timestamp 1666464484
transform 1 0 43332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_471
timestamp 1666464484
transform 1 0 44436 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_483
timestamp 1666464484
transform 1 0 45540 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_488
timestamp 1666464484
transform 1 0 46000 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_500
timestamp 1666464484
transform 1 0 47104 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_512
timestamp 1666464484
transform 1 0 48208 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_524
timestamp 1666464484
transform 1 0 49312 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_536
timestamp 1666464484
transform 1 0 50416 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_548
timestamp 1666464484
transform 1 0 51520 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_553
timestamp 1666464484
transform 1 0 51980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_565
timestamp 1666464484
transform 1 0 53084 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_577
timestamp 1666464484
transform 1 0 54188 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1666464484
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1666464484
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_613
timestamp 1666464484
transform 1 0 57500 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_618
timestamp 1666464484
transform 1 0 57960 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_624
timestamp 1666464484
transform 1 0 58512 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1666464484
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1666464484
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1666464484
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1666464484
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_51
timestamp 1666464484
transform 1 0 5796 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_63
timestamp 1666464484
transform 1 0 6900 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_66
timestamp 1666464484
transform 1 0 7176 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_78
timestamp 1666464484
transform 1 0 8280 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_90
timestamp 1666464484
transform 1 0 9384 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_102
timestamp 1666464484
transform 1 0 10488 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_114
timestamp 1666464484
transform 1 0 11592 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_126
timestamp 1666464484
transform 1 0 12696 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_131
timestamp 1666464484
transform 1 0 13156 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_143
timestamp 1666464484
transform 1 0 14260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_155
timestamp 1666464484
transform 1 0 15364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_167
timestamp 1666464484
transform 1 0 16468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_179
timestamp 1666464484
transform 1 0 17572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_191
timestamp 1666464484
transform 1 0 18676 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_196
timestamp 1666464484
transform 1 0 19136 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_208
timestamp 1666464484
transform 1 0 20240 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_220
timestamp 1666464484
transform 1 0 21344 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_232
timestamp 1666464484
transform 1 0 22448 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_244
timestamp 1666464484
transform 1 0 23552 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_256
timestamp 1666464484
transform 1 0 24656 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1666464484
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_273
timestamp 1666464484
transform 1 0 26220 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_285
timestamp 1666464484
transform 1 0 27324 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_297
timestamp 1666464484
transform 1 0 28428 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_309
timestamp 1666464484
transform 1 0 29532 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_321
timestamp 1666464484
transform 1 0 30636 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_326
timestamp 1666464484
transform 1 0 31096 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_338
timestamp 1666464484
transform 1 0 32200 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_350
timestamp 1666464484
transform 1 0 33304 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_91_379
timestamp 1666464484
transform 1 0 35972 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_387
timestamp 1666464484
transform 1 0 36708 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_391
timestamp 1666464484
transform 1 0 37076 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_403
timestamp 1666464484
transform 1 0 38180 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_415
timestamp 1666464484
transform 1 0 39284 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_427
timestamp 1666464484
transform 1 0 40388 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_439
timestamp 1666464484
transform 1 0 41492 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_451
timestamp 1666464484
transform 1 0 42596 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_456
timestamp 1666464484
transform 1 0 43056 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_468
timestamp 1666464484
transform 1 0 44160 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_480
timestamp 1666464484
transform 1 0 45264 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_492
timestamp 1666464484
transform 1 0 46368 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_504
timestamp 1666464484
transform 1 0 47472 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_516
timestamp 1666464484
transform 1 0 48576 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_521
timestamp 1666464484
transform 1 0 49036 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_533
timestamp 1666464484
transform 1 0 50140 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_545
timestamp 1666464484
transform 1 0 51244 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_557
timestamp 1666464484
transform 1 0 52348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_569
timestamp 1666464484
transform 1 0 53452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_581
timestamp 1666464484
transform 1 0 54556 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_586
timestamp 1666464484
transform 1 0 55016 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_598
timestamp 1666464484
transform 1 0 56120 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_610
timestamp 1666464484
transform 1 0 57224 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_622
timestamp 1666464484
transform 1 0 58328 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1666464484
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1666464484
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_27
timestamp 1666464484
transform 1 0 3588 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_31
timestamp 1666464484
transform 1 0 3956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_33
timestamp 1666464484
transform 1 0 4140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_45
timestamp 1666464484
transform 1 0 5244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_57
timestamp 1666464484
transform 1 0 6348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_69
timestamp 1666464484
transform 1 0 7452 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_81
timestamp 1666464484
transform 1 0 8556 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_93
timestamp 1666464484
transform 1 0 9660 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_98
timestamp 1666464484
transform 1 0 10120 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_110
timestamp 1666464484
transform 1 0 11224 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_122
timestamp 1666464484
transform 1 0 12328 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_134
timestamp 1666464484
transform 1 0 13432 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_146
timestamp 1666464484
transform 1 0 14536 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_158
timestamp 1666464484
transform 1 0 15640 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_163
timestamp 1666464484
transform 1 0 16100 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_175
timestamp 1666464484
transform 1 0 17204 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_187
timestamp 1666464484
transform 1 0 18308 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_199
timestamp 1666464484
transform 1 0 19412 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_211
timestamp 1666464484
transform 1 0 20516 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_223
timestamp 1666464484
transform 1 0 21620 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_228
timestamp 1666464484
transform 1 0 22080 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_240
timestamp 1666464484
transform 1 0 23184 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_252
timestamp 1666464484
transform 1 0 24288 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_264
timestamp 1666464484
transform 1 0 25392 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_276
timestamp 1666464484
transform 1 0 26496 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_288
timestamp 1666464484
transform 1 0 27600 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_293
timestamp 1666464484
transform 1 0 28060 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_305
timestamp 1666464484
transform 1 0 29164 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_317
timestamp 1666464484
transform 1 0 30268 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_329
timestamp 1666464484
transform 1 0 31372 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_341
timestamp 1666464484
transform 1 0 32476 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_353
timestamp 1666464484
transform 1 0 33580 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_358
timestamp 1666464484
transform 1 0 34040 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_370
timestamp 1666464484
transform 1 0 35144 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_382
timestamp 1666464484
transform 1 0 36248 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_394
timestamp 1666464484
transform 1 0 37352 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_406
timestamp 1666464484
transform 1 0 38456 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_418
timestamp 1666464484
transform 1 0 39560 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_423
timestamp 1666464484
transform 1 0 40020 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_435
timestamp 1666464484
transform 1 0 41124 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_447
timestamp 1666464484
transform 1 0 42228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_459
timestamp 1666464484
transform 1 0 43332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_471
timestamp 1666464484
transform 1 0 44436 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_483
timestamp 1666464484
transform 1 0 45540 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_488
timestamp 1666464484
transform 1 0 46000 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_500
timestamp 1666464484
transform 1 0 47104 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_512
timestamp 1666464484
transform 1 0 48208 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_524
timestamp 1666464484
transform 1 0 49312 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_536
timestamp 1666464484
transform 1 0 50416 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_548
timestamp 1666464484
transform 1 0 51520 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_553
timestamp 1666464484
transform 1 0 51980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_565
timestamp 1666464484
transform 1 0 53084 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_577
timestamp 1666464484
transform 1 0 54188 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1666464484
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1666464484
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_613
timestamp 1666464484
transform 1 0 57500 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_92_618
timestamp 1666464484
transform 1 0 57960 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_624
timestamp 1666464484
transform 1 0 58512 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1666464484
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1666464484
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1666464484
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1666464484
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_51
timestamp 1666464484
transform 1 0 5796 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_63
timestamp 1666464484
transform 1 0 6900 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_66
timestamp 1666464484
transform 1 0 7176 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_78
timestamp 1666464484
transform 1 0 8280 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_90
timestamp 1666464484
transform 1 0 9384 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_102
timestamp 1666464484
transform 1 0 10488 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_114
timestamp 1666464484
transform 1 0 11592 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_126
timestamp 1666464484
transform 1 0 12696 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_131
timestamp 1666464484
transform 1 0 13156 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_143
timestamp 1666464484
transform 1 0 14260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_155
timestamp 1666464484
transform 1 0 15364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_167
timestamp 1666464484
transform 1 0 16468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_179
timestamp 1666464484
transform 1 0 17572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_191
timestamp 1666464484
transform 1 0 18676 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_196
timestamp 1666464484
transform 1 0 19136 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_208
timestamp 1666464484
transform 1 0 20240 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_220
timestamp 1666464484
transform 1 0 21344 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_232
timestamp 1666464484
transform 1 0 22448 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_244
timestamp 1666464484
transform 1 0 23552 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_256
timestamp 1666464484
transform 1 0 24656 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1666464484
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_273
timestamp 1666464484
transform 1 0 26220 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_285
timestamp 1666464484
transform 1 0 27324 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_297
timestamp 1666464484
transform 1 0 28428 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_309
timestamp 1666464484
transform 1 0 29532 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_321
timestamp 1666464484
transform 1 0 30636 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_326
timestamp 1666464484
transform 1 0 31096 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_338
timestamp 1666464484
transform 1 0 32200 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_343
timestamp 1666464484
transform 1 0 32660 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_347
timestamp 1666464484
transform 1 0 33028 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_350
timestamp 1666464484
transform 1 0 33304 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_356
timestamp 1666464484
transform 1 0 33856 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_362
timestamp 1666464484
transform 1 0 34408 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_368
timestamp 1666464484
transform 1 0 34960 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_374
timestamp 1666464484
transform 1 0 35512 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_386
timestamp 1666464484
transform 1 0 36616 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_391
timestamp 1666464484
transform 1 0 37076 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_403
timestamp 1666464484
transform 1 0 38180 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_415
timestamp 1666464484
transform 1 0 39284 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_427
timestamp 1666464484
transform 1 0 40388 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_432
timestamp 1666464484
transform 1 0 40848 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_444
timestamp 1666464484
transform 1 0 41952 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_452
timestamp 1666464484
transform 1 0 42688 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_456
timestamp 1666464484
transform 1 0 43056 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_468
timestamp 1666464484
transform 1 0 44160 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_480
timestamp 1666464484
transform 1 0 45264 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_492
timestamp 1666464484
transform 1 0 46368 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_504
timestamp 1666464484
transform 1 0 47472 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_516
timestamp 1666464484
transform 1 0 48576 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_521
timestamp 1666464484
transform 1 0 49036 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_533
timestamp 1666464484
transform 1 0 50140 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_545
timestamp 1666464484
transform 1 0 51244 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_557
timestamp 1666464484
transform 1 0 52348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_569
timestamp 1666464484
transform 1 0 53452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_581
timestamp 1666464484
transform 1 0 54556 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_586
timestamp 1666464484
transform 1 0 55016 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_598
timestamp 1666464484
transform 1 0 56120 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_610
timestamp 1666464484
transform 1 0 57224 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_622
timestamp 1666464484
transform 1 0 58328 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1666464484
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1666464484
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_27
timestamp 1666464484
transform 1 0 3588 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_31
timestamp 1666464484
transform 1 0 3956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_33
timestamp 1666464484
transform 1 0 4140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_45
timestamp 1666464484
transform 1 0 5244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_57
timestamp 1666464484
transform 1 0 6348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_69
timestamp 1666464484
transform 1 0 7452 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_81
timestamp 1666464484
transform 1 0 8556 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_93
timestamp 1666464484
transform 1 0 9660 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_98
timestamp 1666464484
transform 1 0 10120 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_110
timestamp 1666464484
transform 1 0 11224 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_122
timestamp 1666464484
transform 1 0 12328 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_134
timestamp 1666464484
transform 1 0 13432 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_146
timestamp 1666464484
transform 1 0 14536 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_158
timestamp 1666464484
transform 1 0 15640 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_163
timestamp 1666464484
transform 1 0 16100 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_175
timestamp 1666464484
transform 1 0 17204 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_187
timestamp 1666464484
transform 1 0 18308 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_199
timestamp 1666464484
transform 1 0 19412 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_211
timestamp 1666464484
transform 1 0 20516 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_223
timestamp 1666464484
transform 1 0 21620 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_228
timestamp 1666464484
transform 1 0 22080 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_240
timestamp 1666464484
transform 1 0 23184 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_252
timestamp 1666464484
transform 1 0 24288 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_264
timestamp 1666464484
transform 1 0 25392 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_276
timestamp 1666464484
transform 1 0 26496 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_284
timestamp 1666464484
transform 1 0 27232 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_288
timestamp 1666464484
transform 1 0 27600 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_293
timestamp 1666464484
transform 1 0 28060 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_297
timestamp 1666464484
transform 1 0 28428 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_300
timestamp 1666464484
transform 1 0 28704 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_306
timestamp 1666464484
transform 1 0 29256 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_317
timestamp 1666464484
transform 1 0 30268 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_329
timestamp 1666464484
transform 1 0 31372 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_337
timestamp 1666464484
transform 1 0 32108 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_346
timestamp 1666464484
transform 1 0 32936 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_355
timestamp 1666464484
transform 1 0 33764 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_358
timestamp 1666464484
transform 1 0 34040 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_362
timestamp 1666464484
transform 1 0 34408 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_368
timestamp 1666464484
transform 1 0 34960 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_374
timestamp 1666464484
transform 1 0 35512 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_380
timestamp 1666464484
transform 1 0 36064 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_392
timestamp 1666464484
transform 1 0 37168 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_404
timestamp 1666464484
transform 1 0 38272 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_416
timestamp 1666464484
transform 1 0 39376 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_94_423
timestamp 1666464484
transform 1 0 40020 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_427
timestamp 1666464484
transform 1 0 40388 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_433
timestamp 1666464484
transform 1 0 40940 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_439
timestamp 1666464484
transform 1 0 41492 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_448
timestamp 1666464484
transform 1 0 42320 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_460
timestamp 1666464484
transform 1 0 43424 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_472
timestamp 1666464484
transform 1 0 44528 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_484
timestamp 1666464484
transform 1 0 45632 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_488
timestamp 1666464484
transform 1 0 46000 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_500
timestamp 1666464484
transform 1 0 47104 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_512
timestamp 1666464484
transform 1 0 48208 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_524
timestamp 1666464484
transform 1 0 49312 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_536
timestamp 1666464484
transform 1 0 50416 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_548
timestamp 1666464484
transform 1 0 51520 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_553
timestamp 1666464484
transform 1 0 51980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_565
timestamp 1666464484
transform 1 0 53084 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_577
timestamp 1666464484
transform 1 0 54188 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1666464484
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1666464484
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_613
timestamp 1666464484
transform 1 0 57500 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_618
timestamp 1666464484
transform 1 0 57960 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_624
timestamp 1666464484
transform 1 0 58512 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1666464484
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1666464484
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1666464484
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1666464484
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_51
timestamp 1666464484
transform 1 0 5796 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_63
timestamp 1666464484
transform 1 0 6900 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_66
timestamp 1666464484
transform 1 0 7176 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_78
timestamp 1666464484
transform 1 0 8280 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_90
timestamp 1666464484
transform 1 0 9384 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_102
timestamp 1666464484
transform 1 0 10488 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_114
timestamp 1666464484
transform 1 0 11592 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_126
timestamp 1666464484
transform 1 0 12696 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_131
timestamp 1666464484
transform 1 0 13156 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_143
timestamp 1666464484
transform 1 0 14260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_155
timestamp 1666464484
transform 1 0 15364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_167
timestamp 1666464484
transform 1 0 16468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_179
timestamp 1666464484
transform 1 0 17572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_191
timestamp 1666464484
transform 1 0 18676 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_196
timestamp 1666464484
transform 1 0 19136 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_208
timestamp 1666464484
transform 1 0 20240 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_220
timestamp 1666464484
transform 1 0 21344 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_232
timestamp 1666464484
transform 1 0 22448 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_244
timestamp 1666464484
transform 1 0 23552 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_256
timestamp 1666464484
transform 1 0 24656 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1666464484
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_273
timestamp 1666464484
transform 1 0 26220 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_95_278
timestamp 1666464484
transform 1 0 26680 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_286
timestamp 1666464484
transform 1 0 27416 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_292
timestamp 1666464484
transform 1 0 27968 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_303
timestamp 1666464484
transform 1 0 28980 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_312
timestamp 1666464484
transform 1 0 29808 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_323
timestamp 1666464484
transform 1 0 30820 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_326
timestamp 1666464484
transform 1 0 31096 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_330
timestamp 1666464484
transform 1 0 31464 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_95_345
timestamp 1666464484
transform 1 0 32844 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_95_361
timestamp 1666464484
transform 1 0 34316 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_372
timestamp 1666464484
transform 1 0 35328 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_382
timestamp 1666464484
transform 1 0 36248 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_388
timestamp 1666464484
transform 1 0 36800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_391
timestamp 1666464484
transform 1 0 37076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_395
timestamp 1666464484
transform 1 0 37444 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_403
timestamp 1666464484
transform 1 0 38180 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_407
timestamp 1666464484
transform 1 0 38548 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_414
timestamp 1666464484
transform 1 0 39192 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_420
timestamp 1666464484
transform 1 0 39744 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_427
timestamp 1666464484
transform 1 0 40388 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_440
timestamp 1666464484
transform 1 0 41584 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_450
timestamp 1666464484
transform 1 0 42504 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_454
timestamp 1666464484
transform 1 0 42872 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_456
timestamp 1666464484
transform 1 0 43056 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_464
timestamp 1666464484
transform 1 0 43792 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_476
timestamp 1666464484
transform 1 0 44896 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_488
timestamp 1666464484
transform 1 0 46000 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_500
timestamp 1666464484
transform 1 0 47104 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_512
timestamp 1666464484
transform 1 0 48208 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_95_521
timestamp 1666464484
transform 1 0 49036 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_533
timestamp 1666464484
transform 1 0 50140 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_545
timestamp 1666464484
transform 1 0 51244 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_557
timestamp 1666464484
transform 1 0 52348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_569
timestamp 1666464484
transform 1 0 53452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_581
timestamp 1666464484
transform 1 0 54556 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_586
timestamp 1666464484
transform 1 0 55016 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_598
timestamp 1666464484
transform 1 0 56120 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_610
timestamp 1666464484
transform 1 0 57224 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_622
timestamp 1666464484
transform 1 0 58328 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1666464484
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1666464484
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_27
timestamp 1666464484
transform 1 0 3588 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_31
timestamp 1666464484
transform 1 0 3956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_33
timestamp 1666464484
transform 1 0 4140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_45
timestamp 1666464484
transform 1 0 5244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_57
timestamp 1666464484
transform 1 0 6348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_69
timestamp 1666464484
transform 1 0 7452 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_81
timestamp 1666464484
transform 1 0 8556 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_93
timestamp 1666464484
transform 1 0 9660 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_98
timestamp 1666464484
transform 1 0 10120 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_110
timestamp 1666464484
transform 1 0 11224 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_122
timestamp 1666464484
transform 1 0 12328 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_134
timestamp 1666464484
transform 1 0 13432 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_146
timestamp 1666464484
transform 1 0 14536 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_158
timestamp 1666464484
transform 1 0 15640 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_163
timestamp 1666464484
transform 1 0 16100 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_175
timestamp 1666464484
transform 1 0 17204 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_187
timestamp 1666464484
transform 1 0 18308 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_199
timestamp 1666464484
transform 1 0 19412 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_211
timestamp 1666464484
transform 1 0 20516 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_223
timestamp 1666464484
transform 1 0 21620 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_228
timestamp 1666464484
transform 1 0 22080 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_240
timestamp 1666464484
transform 1 0 23184 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_254
timestamp 1666464484
transform 1 0 24472 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_260
timestamp 1666464484
transform 1 0 25024 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_263
timestamp 1666464484
transform 1 0 25300 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_269
timestamp 1666464484
transform 1 0 25852 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_275
timestamp 1666464484
transform 1 0 26404 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_282
timestamp 1666464484
transform 1 0 27048 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_286
timestamp 1666464484
transform 1 0 27416 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_290
timestamp 1666464484
transform 1 0 27784 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_96_293
timestamp 1666464484
transform 1 0 28060 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_300
timestamp 1666464484
transform 1 0 28704 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_311
timestamp 1666464484
transform 1 0 29716 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_318
timestamp 1666464484
transform 1 0 30360 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_326
timestamp 1666464484
transform 1 0 31096 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_334
timestamp 1666464484
transform 1 0 31832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_341
timestamp 1666464484
transform 1 0 32476 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_351
timestamp 1666464484
transform 1 0 33396 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_96_358
timestamp 1666464484
transform 1 0 34040 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_366
timestamp 1666464484
transform 1 0 34776 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_373
timestamp 1666464484
transform 1 0 35420 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_380
timestamp 1666464484
transform 1 0 36064 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_387
timestamp 1666464484
transform 1 0 36708 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_393
timestamp 1666464484
transform 1 0 37260 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_96_402
timestamp 1666464484
transform 1 0 38088 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_408
timestamp 1666464484
transform 1 0 38640 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_96_419
timestamp 1666464484
transform 1 0 39652 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_423
timestamp 1666464484
transform 1 0 40020 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_427
timestamp 1666464484
transform 1 0 40388 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_437
timestamp 1666464484
transform 1 0 41308 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_444
timestamp 1666464484
transform 1 0 41952 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_448
timestamp 1666464484
transform 1 0 42320 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_457
timestamp 1666464484
transform 1 0 43148 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_468
timestamp 1666464484
transform 1 0 44160 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_478
timestamp 1666464484
transform 1 0 45080 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_486
timestamp 1666464484
transform 1 0 45816 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_488
timestamp 1666464484
transform 1 0 46000 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_500
timestamp 1666464484
transform 1 0 47104 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_512
timestamp 1666464484
transform 1 0 48208 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_524
timestamp 1666464484
transform 1 0 49312 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_536
timestamp 1666464484
transform 1 0 50416 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_548
timestamp 1666464484
transform 1 0 51520 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_553
timestamp 1666464484
transform 1 0 51980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_565
timestamp 1666464484
transform 1 0 53084 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_577
timestamp 1666464484
transform 1 0 54188 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1666464484
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1666464484
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_613
timestamp 1666464484
transform 1 0 57500 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_618
timestamp 1666464484
transform 1 0 57960 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_624
timestamp 1666464484
transform 1 0 58512 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1666464484
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1666464484
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1666464484
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1666464484
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_51
timestamp 1666464484
transform 1 0 5796 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_63
timestamp 1666464484
transform 1 0 6900 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_66
timestamp 1666464484
transform 1 0 7176 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_78
timestamp 1666464484
transform 1 0 8280 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_90
timestamp 1666464484
transform 1 0 9384 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_102
timestamp 1666464484
transform 1 0 10488 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_114
timestamp 1666464484
transform 1 0 11592 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_126
timestamp 1666464484
transform 1 0 12696 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_131
timestamp 1666464484
transform 1 0 13156 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_143
timestamp 1666464484
transform 1 0 14260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_155
timestamp 1666464484
transform 1 0 15364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_167
timestamp 1666464484
transform 1 0 16468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_179
timestamp 1666464484
transform 1 0 17572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_191
timestamp 1666464484
transform 1 0 18676 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_196
timestamp 1666464484
transform 1 0 19136 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_208
timestamp 1666464484
transform 1 0 20240 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_220
timestamp 1666464484
transform 1 0 21344 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_232
timestamp 1666464484
transform 1 0 22448 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_244
timestamp 1666464484
transform 1 0 23552 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_97_250
timestamp 1666464484
transform 1 0 24104 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_97_258
timestamp 1666464484
transform 1 0 24840 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_261
timestamp 1666464484
transform 1 0 25116 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_268
timestamp 1666464484
transform 1 0 25760 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_272
timestamp 1666464484
transform 1 0 26128 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_276
timestamp 1666464484
transform 1 0 26496 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_283
timestamp 1666464484
transform 1 0 27140 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_97_291
timestamp 1666464484
transform 1 0 27876 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_297
timestamp 1666464484
transform 1 0 28428 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_304
timestamp 1666464484
transform 1 0 29072 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_308
timestamp 1666464484
transform 1 0 29440 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_314
timestamp 1666464484
transform 1 0 29992 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_323
timestamp 1666464484
transform 1 0 30820 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_97_326
timestamp 1666464484
transform 1 0 31096 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_332
timestamp 1666464484
transform 1 0 31648 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_339
timestamp 1666464484
transform 1 0 32292 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_348
timestamp 1666464484
transform 1 0 33120 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_355
timestamp 1666464484
transform 1 0 33764 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_359
timestamp 1666464484
transform 1 0 34132 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_364
timestamp 1666464484
transform 1 0 34592 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_375
timestamp 1666464484
transform 1 0 35604 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_97_384
timestamp 1666464484
transform 1 0 36432 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_97_391
timestamp 1666464484
transform 1 0 37076 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_97_396
timestamp 1666464484
transform 1 0 37536 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_97_408
timestamp 1666464484
transform 1 0 38640 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_417
timestamp 1666464484
transform 1 0 39468 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_425
timestamp 1666464484
transform 1 0 40204 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_429
timestamp 1666464484
transform 1 0 40572 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_436
timestamp 1666464484
transform 1 0 41216 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_446
timestamp 1666464484
transform 1 0 42136 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_453
timestamp 1666464484
transform 1 0 42780 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_456
timestamp 1666464484
transform 1 0 43056 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_461
timestamp 1666464484
transform 1 0 43516 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_467
timestamp 1666464484
transform 1 0 44068 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_473
timestamp 1666464484
transform 1 0 44620 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_479
timestamp 1666464484
transform 1 0 45172 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1666464484
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_497
timestamp 1666464484
transform 1 0 46828 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_509
timestamp 1666464484
transform 1 0 47932 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_517
timestamp 1666464484
transform 1 0 48668 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_521
timestamp 1666464484
transform 1 0 49036 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_533
timestamp 1666464484
transform 1 0 50140 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_545
timestamp 1666464484
transform 1 0 51244 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_557
timestamp 1666464484
transform 1 0 52348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_569
timestamp 1666464484
transform 1 0 53452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_581
timestamp 1666464484
transform 1 0 54556 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_586
timestamp 1666464484
transform 1 0 55016 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_598
timestamp 1666464484
transform 1 0 56120 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_610
timestamp 1666464484
transform 1 0 57224 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_622
timestamp 1666464484
transform 1 0 58328 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1666464484
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1666464484
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_27
timestamp 1666464484
transform 1 0 3588 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_31
timestamp 1666464484
transform 1 0 3956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_33
timestamp 1666464484
transform 1 0 4140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_45
timestamp 1666464484
transform 1 0 5244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_57
timestamp 1666464484
transform 1 0 6348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_69
timestamp 1666464484
transform 1 0 7452 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_81
timestamp 1666464484
transform 1 0 8556 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_93
timestamp 1666464484
transform 1 0 9660 0 1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_98
timestamp 1666464484
transform 1 0 10120 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_110
timestamp 1666464484
transform 1 0 11224 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_122
timestamp 1666464484
transform 1 0 12328 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_134
timestamp 1666464484
transform 1 0 13432 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_146
timestamp 1666464484
transform 1 0 14536 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_158
timestamp 1666464484
transform 1 0 15640 0 1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_163
timestamp 1666464484
transform 1 0 16100 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_175
timestamp 1666464484
transform 1 0 17204 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_187
timestamp 1666464484
transform 1 0 18308 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_199
timestamp 1666464484
transform 1 0 19412 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_211
timestamp 1666464484
transform 1 0 20516 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_223
timestamp 1666464484
transform 1 0 21620 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_228
timestamp 1666464484
transform 1 0 22080 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_236
timestamp 1666464484
transform 1 0 22816 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_241
timestamp 1666464484
transform 1 0 23276 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_250
timestamp 1666464484
transform 1 0 24104 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_254
timestamp 1666464484
transform 1 0 24472 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_258
timestamp 1666464484
transform 1 0 24840 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_267
timestamp 1666464484
transform 1 0 25668 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_274
timestamp 1666464484
transform 1 0 26312 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_283
timestamp 1666464484
transform 1 0 27140 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_290
timestamp 1666464484
transform 1 0 27784 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_293
timestamp 1666464484
transform 1 0 28060 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_304
timestamp 1666464484
transform 1 0 29072 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_313
timestamp 1666464484
transform 1 0 29900 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_319
timestamp 1666464484
transform 1 0 30452 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_331
timestamp 1666464484
transform 1 0 31556 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_341
timestamp 1666464484
transform 1 0 32476 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_351
timestamp 1666464484
transform 1 0 33396 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_98_358
timestamp 1666464484
transform 1 0 34040 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_364
timestamp 1666464484
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_372
timestamp 1666464484
transform 1 0 35328 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_379
timestamp 1666464484
transform 1 0 35972 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_390
timestamp 1666464484
transform 1 0 36984 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_398
timestamp 1666464484
transform 1 0 37720 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_409
timestamp 1666464484
transform 1 0 38732 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_418
timestamp 1666464484
transform 1 0 39560 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_423
timestamp 1666464484
transform 1 0 40020 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_430
timestamp 1666464484
transform 1 0 40664 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_439
timestamp 1666464484
transform 1 0 41492 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_447
timestamp 1666464484
transform 1 0 42228 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_454
timestamp 1666464484
transform 1 0 42872 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_461
timestamp 1666464484
transform 1 0 43516 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_469
timestamp 1666464484
transform 1 0 44252 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_480
timestamp 1666464484
transform 1 0 45264 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_486
timestamp 1666464484
transform 1 0 45816 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_488
timestamp 1666464484
transform 1 0 46000 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_492
timestamp 1666464484
transform 1 0 46368 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_498
timestamp 1666464484
transform 1 0 46920 0 1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_504
timestamp 1666464484
transform 1 0 47472 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_516
timestamp 1666464484
transform 1 0 48576 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_528
timestamp 1666464484
transform 1 0 49680 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_540
timestamp 1666464484
transform 1 0 50784 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_553
timestamp 1666464484
transform 1 0 51980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_565
timestamp 1666464484
transform 1 0 53084 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_577
timestamp 1666464484
transform 1 0 54188 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1666464484
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1666464484
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_613
timestamp 1666464484
transform 1 0 57500 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_618
timestamp 1666464484
transform 1 0 57960 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_624
timestamp 1666464484
transform 1 0 58512 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1666464484
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1666464484
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1666464484
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1666464484
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_51
timestamp 1666464484
transform 1 0 5796 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_63
timestamp 1666464484
transform 1 0 6900 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_66
timestamp 1666464484
transform 1 0 7176 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_78
timestamp 1666464484
transform 1 0 8280 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_90
timestamp 1666464484
transform 1 0 9384 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_102
timestamp 1666464484
transform 1 0 10488 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_114
timestamp 1666464484
transform 1 0 11592 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_126
timestamp 1666464484
transform 1 0 12696 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_131
timestamp 1666464484
transform 1 0 13156 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_143
timestamp 1666464484
transform 1 0 14260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_155
timestamp 1666464484
transform 1 0 15364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_167
timestamp 1666464484
transform 1 0 16468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_179
timestamp 1666464484
transform 1 0 17572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_191
timestamp 1666464484
transform 1 0 18676 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_196
timestamp 1666464484
transform 1 0 19136 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_208
timestamp 1666464484
transform 1 0 20240 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_220
timestamp 1666464484
transform 1 0 21344 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_99_230
timestamp 1666464484
transform 1 0 22264 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_237
timestamp 1666464484
transform 1 0 22908 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_244
timestamp 1666464484
transform 1 0 23552 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_254
timestamp 1666464484
transform 1 0 24472 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_99_261
timestamp 1666464484
transform 1 0 25116 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_268
timestamp 1666464484
transform 1 0 25760 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_272
timestamp 1666464484
transform 1 0 26128 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_281
timestamp 1666464484
transform 1 0 26956 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_288
timestamp 1666464484
transform 1 0 27600 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_297
timestamp 1666464484
transform 1 0 28428 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_301
timestamp 1666464484
transform 1 0 28796 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_310
timestamp 1666464484
transform 1 0 29624 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_317
timestamp 1666464484
transform 1 0 30268 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_323
timestamp 1666464484
transform 1 0 30820 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_326
timestamp 1666464484
transform 1 0 31096 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_336
timestamp 1666464484
transform 1 0 32016 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_343
timestamp 1666464484
transform 1 0 32660 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_347
timestamp 1666464484
transform 1 0 33028 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_355
timestamp 1666464484
transform 1 0 33764 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_365
timestamp 1666464484
transform 1 0 34684 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_371
timestamp 1666464484
transform 1 0 35236 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_377
timestamp 1666464484
transform 1 0 35788 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_381
timestamp 1666464484
transform 1 0 36156 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_388
timestamp 1666464484
transform 1 0 36800 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_99_391
timestamp 1666464484
transform 1 0 37076 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_99_403
timestamp 1666464484
transform 1 0 38180 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_412
timestamp 1666464484
transform 1 0 39008 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_420
timestamp 1666464484
transform 1 0 39744 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_429
timestamp 1666464484
transform 1 0 40572 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_433
timestamp 1666464484
transform 1 0 40940 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_440
timestamp 1666464484
transform 1 0 41584 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_451
timestamp 1666464484
transform 1 0 42596 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_456
timestamp 1666464484
transform 1 0 43056 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_464
timestamp 1666464484
transform 1 0 43792 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_468
timestamp 1666464484
transform 1 0 44160 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_476
timestamp 1666464484
transform 1 0 44896 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_485
timestamp 1666464484
transform 1 0 45724 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_492
timestamp 1666464484
transform 1 0 46368 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_499
timestamp 1666464484
transform 1 0 47012 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_506
timestamp 1666464484
transform 1 0 47656 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_512
timestamp 1666464484
transform 1 0 48208 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_515
timestamp 1666464484
transform 1 0 48484 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_519
timestamp 1666464484
transform 1 0 48852 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_521
timestamp 1666464484
transform 1 0 49036 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1666464484
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_541
timestamp 1666464484
transform 1 0 50876 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_547
timestamp 1666464484
transform 1 0 51428 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_555
timestamp 1666464484
transform 1 0 52164 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_559
timestamp 1666464484
transform 1 0 52532 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_571
timestamp 1666464484
transform 1 0 53636 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_99_579
timestamp 1666464484
transform 1 0 54372 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_586
timestamp 1666464484
transform 1 0 55016 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_598
timestamp 1666464484
transform 1 0 56120 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_610
timestamp 1666464484
transform 1 0 57224 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_622
timestamp 1666464484
transform 1 0 58328 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1666464484
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1666464484
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_27
timestamp 1666464484
transform 1 0 3588 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_31
timestamp 1666464484
transform 1 0 3956 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_33
timestamp 1666464484
transform 1 0 4140 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_100_42
timestamp 1666464484
transform 1 0 4968 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_50
timestamp 1666464484
transform 1 0 5704 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_62
timestamp 1666464484
transform 1 0 6808 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_74
timestamp 1666464484
transform 1 0 7912 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_86
timestamp 1666464484
transform 1 0 9016 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_94
timestamp 1666464484
transform 1 0 9752 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_100_98
timestamp 1666464484
transform 1 0 10120 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_103
timestamp 1666464484
transform 1 0 10580 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_107
timestamp 1666464484
transform 1 0 10948 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_110
timestamp 1666464484
transform 1 0 11224 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_122
timestamp 1666464484
transform 1 0 12328 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_128
timestamp 1666464484
transform 1 0 12880 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_132
timestamp 1666464484
transform 1 0 13248 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_144
timestamp 1666464484
transform 1 0 14352 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_156
timestamp 1666464484
transform 1 0 15456 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_100_163
timestamp 1666464484
transform 1 0 16100 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_168
timestamp 1666464484
transform 1 0 16560 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_180
timestamp 1666464484
transform 1 0 17664 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_192
timestamp 1666464484
transform 1 0 18768 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_207
timestamp 1666464484
transform 1 0 20148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_222
timestamp 1666464484
transform 1 0 21528 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_226
timestamp 1666464484
transform 1 0 21896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_228
timestamp 1666464484
transform 1 0 22080 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_234
timestamp 1666464484
transform 1 0 22632 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_238
timestamp 1666464484
transform 1 0 23000 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_250
timestamp 1666464484
transform 1 0 24104 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_256
timestamp 1666464484
transform 1 0 24656 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_268
timestamp 1666464484
transform 1 0 25760 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_272
timestamp 1666464484
transform 1 0 26128 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_278
timestamp 1666464484
transform 1 0 26680 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_282
timestamp 1666464484
transform 1 0 27048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_290
timestamp 1666464484
transform 1 0 27784 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_100_293
timestamp 1666464484
transform 1 0 28060 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_300
timestamp 1666464484
transform 1 0 28704 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_313
timestamp 1666464484
transform 1 0 29900 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_321
timestamp 1666464484
transform 1 0 30636 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_329
timestamp 1666464484
transform 1 0 31372 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_341
timestamp 1666464484
transform 1 0 32476 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_351
timestamp 1666464484
transform 1 0 33396 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_100_358
timestamp 1666464484
transform 1 0 34040 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_363
timestamp 1666464484
transform 1 0 34500 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_375
timestamp 1666464484
transform 1 0 35604 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_389
timestamp 1666464484
transform 1 0 36892 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_397
timestamp 1666464484
transform 1 0 37628 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_405
timestamp 1666464484
transform 1 0 38364 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_100_419
timestamp 1666464484
transform 1 0 39652 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_100_423
timestamp 1666464484
transform 1 0 40020 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_431
timestamp 1666464484
transform 1 0 40756 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_443
timestamp 1666464484
transform 1 0 41860 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_449
timestamp 1666464484
transform 1 0 42412 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_459
timestamp 1666464484
transform 1 0 43332 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_473
timestamp 1666464484
transform 1 0 44620 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_480
timestamp 1666464484
transform 1 0 45264 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_486
timestamp 1666464484
transform 1 0 45816 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_488
timestamp 1666464484
transform 1 0 46000 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_493
timestamp 1666464484
transform 1 0 46460 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_500
timestamp 1666464484
transform 1 0 47104 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_507
timestamp 1666464484
transform 1 0 47748 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_514
timestamp 1666464484
transform 1 0 48392 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_521
timestamp 1666464484
transform 1 0 49036 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_528
timestamp 1666464484
transform 1 0 49680 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_535
timestamp 1666464484
transform 1 0 50324 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_542
timestamp 1666464484
transform 1 0 50968 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_100_549
timestamp 1666464484
transform 1 0 51612 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_100_553
timestamp 1666464484
transform 1 0 51980 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_558
timestamp 1666464484
transform 1 0 52440 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_565
timestamp 1666464484
transform 1 0 53084 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_572
timestamp 1666464484
transform 1 0 53728 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_578
timestamp 1666464484
transform 1 0 54280 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_582
timestamp 1666464484
transform 1 0 54648 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_589
timestamp 1666464484
transform 1 0 55292 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_595
timestamp 1666464484
transform 1 0 55844 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_602
timestamp 1666464484
transform 1 0 56488 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_614
timestamp 1666464484
transform 1 0 57592 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_100_618
timestamp 1666464484
transform 1 0 57960 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_624
timestamp 1666464484
transform 1 0 58512 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1666464484
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1666464484
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 1666464484
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_30
timestamp 1666464484
transform 1 0 3864 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_33
timestamp 1666464484
transform 1 0 4140 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_39
timestamp 1666464484
transform 1 0 4692 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_43
timestamp 1666464484
transform 1 0 5060 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_48
timestamp 1666464484
transform 1 0 5520 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_55
timestamp 1666464484
transform 1 0 6164 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_62
timestamp 1666464484
transform 1 0 6808 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_65
timestamp 1666464484
transform 1 0 7084 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_70
timestamp 1666464484
transform 1 0 7544 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_77
timestamp 1666464484
transform 1 0 8188 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_81
timestamp 1666464484
transform 1 0 8556 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_85
timestamp 1666464484
transform 1 0 8924 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_92
timestamp 1666464484
transform 1 0 9568 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_97
timestamp 1666464484
transform 1 0 10028 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_103
timestamp 1666464484
transform 1 0 10580 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_108
timestamp 1666464484
transform 1 0 11040 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_115
timestamp 1666464484
transform 1 0 11684 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_123
timestamp 1666464484
transform 1 0 12420 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_127
timestamp 1666464484
transform 1 0 12788 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_129
timestamp 1666464484
transform 1 0 12972 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_133
timestamp 1666464484
transform 1 0 13340 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_138
timestamp 1666464484
transform 1 0 13800 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_145
timestamp 1666464484
transform 1 0 14444 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_153
timestamp 1666464484
transform 1 0 15180 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_159
timestamp 1666464484
transform 1 0 15732 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_161
timestamp 1666464484
transform 1 0 15916 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_168
timestamp 1666464484
transform 1 0 16560 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_175
timestamp 1666464484
transform 1 0 17204 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_183
timestamp 1666464484
transform 1 0 17940 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_190
timestamp 1666464484
transform 1 0 18584 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_193
timestamp 1666464484
transform 1 0 18860 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_199
timestamp 1666464484
transform 1 0 19412 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_207
timestamp 1666464484
transform 1 0 20148 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_213
timestamp 1666464484
transform 1 0 20700 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_101_222
timestamp 1666464484
transform 1 0 21528 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_225
timestamp 1666464484
transform 1 0 21804 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_231
timestamp 1666464484
transform 1 0 22356 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_243
timestamp 1666464484
transform 1 0 23460 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_252
timestamp 1666464484
transform 1 0 24288 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_257
timestamp 1666464484
transform 1 0 24748 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_263
timestamp 1666464484
transform 1 0 25300 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_273
timestamp 1666464484
transform 1 0 26220 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_279
timestamp 1666464484
transform 1 0 26772 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_286
timestamp 1666464484
transform 1 0 27416 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_289
timestamp 1666464484
transform 1 0 27692 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_295
timestamp 1666464484
transform 1 0 28244 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_303
timestamp 1666464484
transform 1 0 28980 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_307
timestamp 1666464484
transform 1 0 29348 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_311
timestamp 1666464484
transform 1 0 29716 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_318
timestamp 1666464484
transform 1 0 30360 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_101_321
timestamp 1666464484
transform 1 0 30636 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_327
timestamp 1666464484
transform 1 0 31188 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_333
timestamp 1666464484
transform 1 0 31740 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_344
timestamp 1666464484
transform 1 0 32752 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_350
timestamp 1666464484
transform 1 0 33304 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_353
timestamp 1666464484
transform 1 0 33580 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_361
timestamp 1666464484
transform 1 0 34316 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_369
timestamp 1666464484
transform 1 0 35052 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_376
timestamp 1666464484
transform 1 0 35696 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_382
timestamp 1666464484
transform 1 0 36248 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_385
timestamp 1666464484
transform 1 0 36524 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_397
timestamp 1666464484
transform 1 0 37628 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_411
timestamp 1666464484
transform 1 0 38916 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_415
timestamp 1666464484
transform 1 0 39284 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_417
timestamp 1666464484
transform 1 0 39468 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_430
timestamp 1666464484
transform 1 0 40664 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_437
timestamp 1666464484
transform 1 0 41308 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_446
timestamp 1666464484
transform 1 0 42136 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_449
timestamp 1666464484
transform 1 0 42412 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_453
timestamp 1666464484
transform 1 0 42780 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_464
timestamp 1666464484
transform 1 0 43792 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_471
timestamp 1666464484
transform 1 0 44436 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_478
timestamp 1666464484
transform 1 0 45080 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_101_481
timestamp 1666464484
transform 1 0 45356 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_488
timestamp 1666464484
transform 1 0 46000 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_495
timestamp 1666464484
transform 1 0 46644 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_101_509
timestamp 1666464484
transform 1 0 47932 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_513
timestamp 1666464484
transform 1 0 48300 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_525
timestamp 1666464484
transform 1 0 49404 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_539
timestamp 1666464484
transform 1 0 50692 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_543
timestamp 1666464484
transform 1 0 51060 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_545
timestamp 1666464484
transform 1 0 51244 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_551
timestamp 1666464484
transform 1 0 51796 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_565
timestamp 1666464484
transform 1 0 53084 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_572
timestamp 1666464484
transform 1 0 53728 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_577
timestamp 1666464484
transform 1 0 54188 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_583
timestamp 1666464484
transform 1 0 54740 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_593
timestamp 1666464484
transform 1 0 55660 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_600
timestamp 1666464484
transform 1 0 56304 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_609
timestamp 1666464484
transform 1 0 57132 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_621
timestamp 1666464484
transform 1 0 58236 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666464484
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666464484
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666464484
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666464484
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666464484
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666464484
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666464484
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666464484
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666464484
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666464484
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666464484
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666464484
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666464484
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666464484
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666464484
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666464484
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666464484
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666464484
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666464484
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666464484
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666464484
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666464484
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666464484
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666464484
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666464484
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666464484
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666464484
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666464484
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666464484
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666464484
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666464484
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666464484
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666464484
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666464484
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666464484
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666464484
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1666464484
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1666464484
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1666464484
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1666464484
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1666464484
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1666464484
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1666464484
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1666464484
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1666464484
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1666464484
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1666464484
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1666464484
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1666464484
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1666464484
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1666464484
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1666464484
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1666464484
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1666464484
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1666464484
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1666464484
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1666464484
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1666464484
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1666464484
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1666464484
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1666464484
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1666464484
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1666464484
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1666464484
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1666464484
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1666464484
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1666464484
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1666464484
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1666464484
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1666464484
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1666464484
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1666464484
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1666464484
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1666464484
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 6992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 9936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 12880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 15824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 18768 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 24656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 27600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 30544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 33488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 36432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 39376 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 45264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 48208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 51152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 54096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 57040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 13064 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 19044 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 25024 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 31004 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 36984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 42964 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 48944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 54924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 4048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 16008 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 21988 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 27968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 33948 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 39928 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 45908 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 51888 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 57868 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 13064 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 19044 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 25024 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 31004 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 36984 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 42964 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 48944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 54924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 4048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 16008 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 21988 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 27968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 33948 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 39928 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 45908 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 51888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 57868 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 13064 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 19044 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 25024 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 31004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 36984 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 42964 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 48944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 54924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 4048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 16008 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 21988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 27968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 33948 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 39928 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 45908 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 51888 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 57868 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 13064 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 19044 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 25024 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 31004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 36984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 42964 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 48944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 54924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 4048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 16008 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 21988 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 27968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 33948 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 39928 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 45908 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 51888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 57868 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 13064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 19044 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 25024 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 31004 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 36984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 42964 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 48944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 54924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 4048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 16008 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 21988 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 27968 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 33948 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 39928 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 45908 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 51888 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 57868 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 7084 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 13064 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 19044 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 25024 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 31004 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 36984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 42964 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 48944 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 54924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 4048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 16008 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 21988 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 27968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 33948 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 39928 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 45908 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 51888 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 57868 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 13064 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 19044 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 25024 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 31004 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 36984 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 42964 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 48944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 54924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 4048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 16008 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 21988 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 27968 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 33948 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 39928 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 45908 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 51888 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 57868 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 13064 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 19044 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 25024 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 31004 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 36984 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 42964 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 48944 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 54924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 4048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 16008 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 21988 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 27968 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 33948 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 39928 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 45908 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 51888 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 57868 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 13064 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 19044 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 25024 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 31004 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 36984 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 42964 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 48944 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 54924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 4048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 16008 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 21988 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 27968 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 33948 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 39928 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 45908 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 51888 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 57868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 13064 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 19044 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 25024 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 31004 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 36984 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 42964 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 48944 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 54924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 4048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 16008 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 21988 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 27968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 33948 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 39928 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 45908 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 51888 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 57868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 13064 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 19044 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 25024 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 31004 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 36984 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 42964 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 48944 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 54924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 4048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 16008 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 21988 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 27968 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 33948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 39928 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 45908 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 51888 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 57868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 7084 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 13064 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 19044 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 25024 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 31004 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 36984 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 42964 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 48944 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 54924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 4048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 16008 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 21988 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 27968 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 33948 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 39928 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 45908 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 51888 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 57868 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 13064 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 19044 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 25024 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 31004 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 36984 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 42964 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 48944 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 54924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 4048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 16008 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 21988 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 27968 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 33948 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 39928 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 45908 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 51888 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 57868 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 7084 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 13064 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 19044 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 25024 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 31004 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 36984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 42964 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 48944 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 54924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 4048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 16008 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 21988 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 27968 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 33948 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 39928 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 45908 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 51888 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 57868 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 7084 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 13064 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 19044 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 25024 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 31004 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 36984 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 42964 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 48944 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 54924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 4048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 16008 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 21988 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 27968 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 33948 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 39928 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 45908 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 51888 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 57868 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 7084 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 13064 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 19044 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 25024 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 31004 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 36984 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 42964 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 48944 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 54924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 4048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 16008 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 21988 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 27968 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 33948 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 39928 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 45908 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 51888 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 57868 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 7084 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 13064 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 19044 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 25024 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 31004 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 36984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 42964 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 48944 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 54924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 4048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 16008 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 21988 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 27968 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 33948 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 39928 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 45908 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 51888 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 57868 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 7084 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 13064 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 19044 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 25024 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 31004 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 36984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 42964 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 48944 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 54924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 4048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 16008 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 21988 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 27968 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 33948 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 39928 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 45908 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 51888 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666464484
transform 1 0 57868 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666464484
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666464484
transform 1 0 13064 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666464484
transform 1 0 19044 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666464484
transform 1 0 25024 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666464484
transform 1 0 31004 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666464484
transform 1 0 36984 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666464484
transform 1 0 42964 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666464484
transform 1 0 48944 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666464484
transform 1 0 54924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666464484
transform 1 0 4048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666464484
transform 1 0 16008 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666464484
transform 1 0 21988 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666464484
transform 1 0 27968 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666464484
transform 1 0 33948 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666464484
transform 1 0 39928 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666464484
transform 1 0 45908 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666464484
transform 1 0 51888 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666464484
transform 1 0 57868 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666464484
transform 1 0 7084 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666464484
transform 1 0 13064 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666464484
transform 1 0 19044 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666464484
transform 1 0 25024 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666464484
transform 1 0 31004 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666464484
transform 1 0 36984 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666464484
transform 1 0 42964 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666464484
transform 1 0 48944 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666464484
transform 1 0 54924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666464484
transform 1 0 4048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666464484
transform 1 0 16008 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666464484
transform 1 0 21988 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666464484
transform 1 0 27968 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666464484
transform 1 0 33948 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666464484
transform 1 0 39928 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666464484
transform 1 0 45908 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666464484
transform 1 0 51888 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666464484
transform 1 0 57868 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666464484
transform 1 0 7084 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666464484
transform 1 0 13064 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666464484
transform 1 0 19044 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666464484
transform 1 0 25024 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666464484
transform 1 0 31004 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666464484
transform 1 0 36984 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666464484
transform 1 0 42964 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666464484
transform 1 0 48944 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666464484
transform 1 0 54924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666464484
transform 1 0 4048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666464484
transform 1 0 16008 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666464484
transform 1 0 21988 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666464484
transform 1 0 27968 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666464484
transform 1 0 33948 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666464484
transform 1 0 39928 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666464484
transform 1 0 45908 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666464484
transform 1 0 51888 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666464484
transform 1 0 57868 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666464484
transform 1 0 7084 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666464484
transform 1 0 13064 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666464484
transform 1 0 19044 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666464484
transform 1 0 25024 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666464484
transform 1 0 31004 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666464484
transform 1 0 36984 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666464484
transform 1 0 42964 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666464484
transform 1 0 48944 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666464484
transform 1 0 54924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666464484
transform 1 0 4048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666464484
transform 1 0 10028 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666464484
transform 1 0 16008 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666464484
transform 1 0 21988 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666464484
transform 1 0 27968 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666464484
transform 1 0 33948 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666464484
transform 1 0 39928 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666464484
transform 1 0 45908 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666464484
transform 1 0 51888 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666464484
transform 1 0 57868 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666464484
transform 1 0 7084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666464484
transform 1 0 13064 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666464484
transform 1 0 19044 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666464484
transform 1 0 25024 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666464484
transform 1 0 31004 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666464484
transform 1 0 36984 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666464484
transform 1 0 42964 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666464484
transform 1 0 48944 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666464484
transform 1 0 54924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666464484
transform 1 0 4048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666464484
transform 1 0 10028 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666464484
transform 1 0 16008 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666464484
transform 1 0 21988 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666464484
transform 1 0 27968 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666464484
transform 1 0 33948 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666464484
transform 1 0 39928 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666464484
transform 1 0 45908 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666464484
transform 1 0 51888 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666464484
transform 1 0 57868 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666464484
transform 1 0 7084 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666464484
transform 1 0 13064 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666464484
transform 1 0 19044 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666464484
transform 1 0 25024 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666464484
transform 1 0 31004 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666464484
transform 1 0 36984 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666464484
transform 1 0 42964 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666464484
transform 1 0 48944 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666464484
transform 1 0 54924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666464484
transform 1 0 4048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666464484
transform 1 0 10028 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666464484
transform 1 0 16008 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666464484
transform 1 0 21988 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666464484
transform 1 0 27968 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666464484
transform 1 0 33948 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666464484
transform 1 0 39928 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666464484
transform 1 0 45908 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666464484
transform 1 0 51888 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666464484
transform 1 0 57868 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666464484
transform 1 0 7084 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666464484
transform 1 0 13064 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666464484
transform 1 0 19044 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666464484
transform 1 0 25024 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666464484
transform 1 0 31004 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666464484
transform 1 0 36984 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666464484
transform 1 0 42964 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666464484
transform 1 0 48944 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666464484
transform 1 0 54924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666464484
transform 1 0 4048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666464484
transform 1 0 10028 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666464484
transform 1 0 16008 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666464484
transform 1 0 21988 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666464484
transform 1 0 27968 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666464484
transform 1 0 33948 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666464484
transform 1 0 39928 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666464484
transform 1 0 45908 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666464484
transform 1 0 51888 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666464484
transform 1 0 57868 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666464484
transform 1 0 7084 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666464484
transform 1 0 13064 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666464484
transform 1 0 19044 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666464484
transform 1 0 25024 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666464484
transform 1 0 31004 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666464484
transform 1 0 36984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666464484
transform 1 0 42964 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666464484
transform 1 0 48944 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666464484
transform 1 0 54924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666464484
transform 1 0 4048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666464484
transform 1 0 10028 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666464484
transform 1 0 16008 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666464484
transform 1 0 21988 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666464484
transform 1 0 27968 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666464484
transform 1 0 33948 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666464484
transform 1 0 39928 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666464484
transform 1 0 45908 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666464484
transform 1 0 51888 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666464484
transform 1 0 57868 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666464484
transform 1 0 7084 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666464484
transform 1 0 13064 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666464484
transform 1 0 19044 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666464484
transform 1 0 25024 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666464484
transform 1 0 31004 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666464484
transform 1 0 36984 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666464484
transform 1 0 42964 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666464484
transform 1 0 48944 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666464484
transform 1 0 54924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666464484
transform 1 0 4048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666464484
transform 1 0 10028 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666464484
transform 1 0 16008 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666464484
transform 1 0 21988 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666464484
transform 1 0 27968 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666464484
transform 1 0 33948 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666464484
transform 1 0 39928 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666464484
transform 1 0 45908 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666464484
transform 1 0 51888 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666464484
transform 1 0 57868 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666464484
transform 1 0 7084 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666464484
transform 1 0 13064 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666464484
transform 1 0 19044 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666464484
transform 1 0 25024 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666464484
transform 1 0 31004 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666464484
transform 1 0 36984 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666464484
transform 1 0 42964 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666464484
transform 1 0 48944 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666464484
transform 1 0 54924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666464484
transform 1 0 4048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666464484
transform 1 0 10028 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666464484
transform 1 0 16008 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666464484
transform 1 0 21988 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666464484
transform 1 0 27968 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666464484
transform 1 0 33948 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666464484
transform 1 0 39928 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666464484
transform 1 0 45908 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666464484
transform 1 0 51888 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666464484
transform 1 0 57868 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666464484
transform 1 0 7084 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666464484
transform 1 0 13064 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666464484
transform 1 0 19044 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666464484
transform 1 0 25024 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666464484
transform 1 0 31004 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666464484
transform 1 0 36984 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666464484
transform 1 0 42964 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666464484
transform 1 0 48944 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666464484
transform 1 0 54924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666464484
transform 1 0 4048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666464484
transform 1 0 10028 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666464484
transform 1 0 16008 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666464484
transform 1 0 21988 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666464484
transform 1 0 27968 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666464484
transform 1 0 33948 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666464484
transform 1 0 39928 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666464484
transform 1 0 45908 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666464484
transform 1 0 51888 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666464484
transform 1 0 57868 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666464484
transform 1 0 7084 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666464484
transform 1 0 13064 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666464484
transform 1 0 19044 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666464484
transform 1 0 25024 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666464484
transform 1 0 31004 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666464484
transform 1 0 36984 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666464484
transform 1 0 42964 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666464484
transform 1 0 48944 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666464484
transform 1 0 54924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666464484
transform 1 0 4048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666464484
transform 1 0 10028 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666464484
transform 1 0 16008 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666464484
transform 1 0 21988 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666464484
transform 1 0 27968 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666464484
transform 1 0 33948 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666464484
transform 1 0 39928 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666464484
transform 1 0 45908 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666464484
transform 1 0 51888 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666464484
transform 1 0 57868 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666464484
transform 1 0 7084 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666464484
transform 1 0 13064 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666464484
transform 1 0 19044 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666464484
transform 1 0 25024 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666464484
transform 1 0 31004 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666464484
transform 1 0 36984 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666464484
transform 1 0 42964 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666464484
transform 1 0 48944 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666464484
transform 1 0 54924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666464484
transform 1 0 4048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666464484
transform 1 0 10028 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666464484
transform 1 0 16008 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666464484
transform 1 0 21988 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666464484
transform 1 0 27968 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666464484
transform 1 0 33948 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666464484
transform 1 0 39928 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666464484
transform 1 0 45908 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666464484
transform 1 0 51888 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666464484
transform 1 0 57868 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666464484
transform 1 0 7084 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666464484
transform 1 0 13064 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666464484
transform 1 0 19044 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666464484
transform 1 0 25024 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666464484
transform 1 0 31004 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666464484
transform 1 0 36984 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666464484
transform 1 0 42964 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666464484
transform 1 0 48944 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666464484
transform 1 0 54924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666464484
transform 1 0 4048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666464484
transform 1 0 10028 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666464484
transform 1 0 16008 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666464484
transform 1 0 21988 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666464484
transform 1 0 27968 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666464484
transform 1 0 33948 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666464484
transform 1 0 39928 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666464484
transform 1 0 45908 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666464484
transform 1 0 51888 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666464484
transform 1 0 57868 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666464484
transform 1 0 7084 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666464484
transform 1 0 13064 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666464484
transform 1 0 19044 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666464484
transform 1 0 25024 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666464484
transform 1 0 31004 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666464484
transform 1 0 36984 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666464484
transform 1 0 42964 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666464484
transform 1 0 48944 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666464484
transform 1 0 54924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666464484
transform 1 0 4048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666464484
transform 1 0 10028 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666464484
transform 1 0 16008 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666464484
transform 1 0 21988 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666464484
transform 1 0 27968 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666464484
transform 1 0 33948 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666464484
transform 1 0 39928 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666464484
transform 1 0 45908 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666464484
transform 1 0 51888 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666464484
transform 1 0 57868 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666464484
transform 1 0 7084 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666464484
transform 1 0 13064 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666464484
transform 1 0 19044 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666464484
transform 1 0 25024 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666464484
transform 1 0 31004 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666464484
transform 1 0 36984 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666464484
transform 1 0 42964 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666464484
transform 1 0 48944 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666464484
transform 1 0 54924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666464484
transform 1 0 4048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666464484
transform 1 0 10028 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666464484
transform 1 0 16008 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666464484
transform 1 0 21988 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666464484
transform 1 0 27968 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666464484
transform 1 0 33948 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666464484
transform 1 0 39928 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666464484
transform 1 0 45908 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666464484
transform 1 0 51888 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666464484
transform 1 0 57868 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666464484
transform 1 0 7084 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666464484
transform 1 0 13064 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666464484
transform 1 0 19044 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666464484
transform 1 0 25024 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666464484
transform 1 0 31004 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666464484
transform 1 0 36984 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666464484
transform 1 0 42964 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666464484
transform 1 0 48944 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666464484
transform 1 0 54924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666464484
transform 1 0 4048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666464484
transform 1 0 10028 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666464484
transform 1 0 16008 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666464484
transform 1 0 21988 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666464484
transform 1 0 27968 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666464484
transform 1 0 33948 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666464484
transform 1 0 39928 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666464484
transform 1 0 45908 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666464484
transform 1 0 51888 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666464484
transform 1 0 57868 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666464484
transform 1 0 7084 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666464484
transform 1 0 13064 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666464484
transform 1 0 19044 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666464484
transform 1 0 25024 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666464484
transform 1 0 31004 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666464484
transform 1 0 36984 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666464484
transform 1 0 42964 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666464484
transform 1 0 48944 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666464484
transform 1 0 54924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666464484
transform 1 0 4048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666464484
transform 1 0 10028 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666464484
transform 1 0 16008 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666464484
transform 1 0 21988 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666464484
transform 1 0 27968 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666464484
transform 1 0 33948 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666464484
transform 1 0 39928 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666464484
transform 1 0 45908 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666464484
transform 1 0 51888 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666464484
transform 1 0 57868 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666464484
transform 1 0 7084 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666464484
transform 1 0 13064 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666464484
transform 1 0 19044 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666464484
transform 1 0 25024 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666464484
transform 1 0 31004 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666464484
transform 1 0 36984 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666464484
transform 1 0 42964 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666464484
transform 1 0 48944 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666464484
transform 1 0 54924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666464484
transform 1 0 4048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666464484
transform 1 0 10028 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666464484
transform 1 0 16008 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666464484
transform 1 0 21988 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666464484
transform 1 0 27968 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666464484
transform 1 0 33948 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666464484
transform 1 0 39928 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666464484
transform 1 0 45908 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666464484
transform 1 0 51888 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666464484
transform 1 0 57868 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666464484
transform 1 0 7084 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666464484
transform 1 0 13064 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666464484
transform 1 0 19044 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666464484
transform 1 0 25024 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666464484
transform 1 0 31004 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1666464484
transform 1 0 36984 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1666464484
transform 1 0 42964 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1666464484
transform 1 0 48944 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1666464484
transform 1 0 54924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1666464484
transform 1 0 4048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1666464484
transform 1 0 10028 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1666464484
transform 1 0 16008 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1666464484
transform 1 0 21988 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1666464484
transform 1 0 27968 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1666464484
transform 1 0 33948 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1666464484
transform 1 0 39928 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1666464484
transform 1 0 45908 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1666464484
transform 1 0 51888 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1666464484
transform 1 0 57868 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1666464484
transform 1 0 7084 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1666464484
transform 1 0 13064 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1666464484
transform 1 0 19044 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1666464484
transform 1 0 25024 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1666464484
transform 1 0 31004 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1666464484
transform 1 0 36984 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1666464484
transform 1 0 42964 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1666464484
transform 1 0 48944 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1666464484
transform 1 0 54924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1666464484
transform 1 0 4048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1666464484
transform 1 0 10028 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1666464484
transform 1 0 16008 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1666464484
transform 1 0 21988 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1666464484
transform 1 0 27968 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1666464484
transform 1 0 33948 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1666464484
transform 1 0 39928 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1666464484
transform 1 0 45908 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1666464484
transform 1 0 51888 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1666464484
transform 1 0 57868 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1666464484
transform 1 0 7084 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1666464484
transform 1 0 13064 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1666464484
transform 1 0 19044 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1666464484
transform 1 0 25024 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1666464484
transform 1 0 31004 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1666464484
transform 1 0 36984 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1666464484
transform 1 0 42964 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1666464484
transform 1 0 48944 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1666464484
transform 1 0 54924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1666464484
transform 1 0 4048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1666464484
transform 1 0 10028 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1666464484
transform 1 0 16008 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1666464484
transform 1 0 21988 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1666464484
transform 1 0 27968 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1666464484
transform 1 0 33948 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1666464484
transform 1 0 39928 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1666464484
transform 1 0 45908 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1666464484
transform 1 0 51888 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1666464484
transform 1 0 57868 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1666464484
transform 1 0 7084 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1666464484
transform 1 0 13064 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1666464484
transform 1 0 19044 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1666464484
transform 1 0 25024 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1666464484
transform 1 0 31004 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1666464484
transform 1 0 36984 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1666464484
transform 1 0 42964 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1666464484
transform 1 0 48944 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1666464484
transform 1 0 54924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1666464484
transform 1 0 4048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1666464484
transform 1 0 10028 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1666464484
transform 1 0 16008 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1666464484
transform 1 0 21988 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1666464484
transform 1 0 27968 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1666464484
transform 1 0 33948 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1666464484
transform 1 0 39928 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1666464484
transform 1 0 45908 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1666464484
transform 1 0 51888 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1666464484
transform 1 0 57868 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1666464484
transform 1 0 7084 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1666464484
transform 1 0 13064 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1666464484
transform 1 0 19044 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1666464484
transform 1 0 25024 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1666464484
transform 1 0 31004 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1666464484
transform 1 0 36984 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1666464484
transform 1 0 42964 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1666464484
transform 1 0 48944 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1666464484
transform 1 0 54924 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1666464484
transform 1 0 4048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1666464484
transform 1 0 10028 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1666464484
transform 1 0 16008 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1666464484
transform 1 0 21988 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1666464484
transform 1 0 27968 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1666464484
transform 1 0 33948 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1666464484
transform 1 0 39928 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1666464484
transform 1 0 45908 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1666464484
transform 1 0 51888 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1666464484
transform 1 0 57868 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1666464484
transform 1 0 7084 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1666464484
transform 1 0 13064 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1666464484
transform 1 0 19044 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1666464484
transform 1 0 25024 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1666464484
transform 1 0 31004 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1666464484
transform 1 0 36984 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1666464484
transform 1 0 42964 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1666464484
transform 1 0 48944 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1666464484
transform 1 0 54924 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1666464484
transform 1 0 4048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1666464484
transform 1 0 10028 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1666464484
transform 1 0 16008 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1666464484
transform 1 0 21988 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1666464484
transform 1 0 27968 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1666464484
transform 1 0 33948 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1666464484
transform 1 0 39928 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1666464484
transform 1 0 45908 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1666464484
transform 1 0 51888 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1666464484
transform 1 0 57868 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1666464484
transform 1 0 7084 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1666464484
transform 1 0 13064 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1666464484
transform 1 0 19044 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1666464484
transform 1 0 25024 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1666464484
transform 1 0 31004 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1666464484
transform 1 0 36984 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1666464484
transform 1 0 42964 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1666464484
transform 1 0 48944 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1666464484
transform 1 0 54924 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1666464484
transform 1 0 4048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1666464484
transform 1 0 10028 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1666464484
transform 1 0 16008 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1666464484
transform 1 0 21988 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1666464484
transform 1 0 27968 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1666464484
transform 1 0 33948 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1666464484
transform 1 0 39928 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1666464484
transform 1 0 45908 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1666464484
transform 1 0 51888 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1666464484
transform 1 0 57868 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1666464484
transform 1 0 7084 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1666464484
transform 1 0 13064 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1666464484
transform 1 0 19044 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1666464484
transform 1 0 25024 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1666464484
transform 1 0 31004 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1666464484
transform 1 0 36984 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1666464484
transform 1 0 42964 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1666464484
transform 1 0 48944 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1666464484
transform 1 0 54924 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1666464484
transform 1 0 4048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1666464484
transform 1 0 10028 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1666464484
transform 1 0 16008 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1666464484
transform 1 0 21988 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1666464484
transform 1 0 27968 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1666464484
transform 1 0 33948 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1666464484
transform 1 0 39928 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1666464484
transform 1 0 45908 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1666464484
transform 1 0 51888 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1666464484
transform 1 0 57868 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1666464484
transform 1 0 7084 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1666464484
transform 1 0 13064 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1666464484
transform 1 0 19044 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1666464484
transform 1 0 25024 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1666464484
transform 1 0 31004 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1666464484
transform 1 0 36984 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1666464484
transform 1 0 42964 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1666464484
transform 1 0 48944 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1666464484
transform 1 0 54924 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1666464484
transform 1 0 4048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1666464484
transform 1 0 10028 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1666464484
transform 1 0 16008 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1666464484
transform 1 0 21988 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1666464484
transform 1 0 27968 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1666464484
transform 1 0 33948 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1666464484
transform 1 0 39928 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1666464484
transform 1 0 45908 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1666464484
transform 1 0 51888 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1666464484
transform 1 0 57868 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1666464484
transform 1 0 7084 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1666464484
transform 1 0 13064 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1666464484
transform 1 0 19044 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1666464484
transform 1 0 25024 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1666464484
transform 1 0 31004 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1666464484
transform 1 0 36984 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1666464484
transform 1 0 42964 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1666464484
transform 1 0 48944 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1666464484
transform 1 0 54924 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1666464484
transform 1 0 4048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1666464484
transform 1 0 10028 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1666464484
transform 1 0 16008 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1666464484
transform 1 0 21988 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1666464484
transform 1 0 27968 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1666464484
transform 1 0 33948 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1666464484
transform 1 0 39928 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1666464484
transform 1 0 45908 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1666464484
transform 1 0 51888 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1666464484
transform 1 0 57868 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1666464484
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1666464484
transform 1 0 13064 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1666464484
transform 1 0 19044 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1666464484
transform 1 0 25024 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1666464484
transform 1 0 31004 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1666464484
transform 1 0 36984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1666464484
transform 1 0 42964 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1666464484
transform 1 0 48944 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1666464484
transform 1 0 54924 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1666464484
transform 1 0 4048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1666464484
transform 1 0 10028 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1666464484
transform 1 0 16008 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1666464484
transform 1 0 21988 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1666464484
transform 1 0 27968 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1666464484
transform 1 0 33948 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1666464484
transform 1 0 39928 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1666464484
transform 1 0 45908 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1666464484
transform 1 0 51888 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1666464484
transform 1 0 57868 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1666464484
transform 1 0 7084 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1666464484
transform 1 0 13064 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1666464484
transform 1 0 19044 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1666464484
transform 1 0 25024 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1666464484
transform 1 0 31004 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1666464484
transform 1 0 36984 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1666464484
transform 1 0 42964 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1666464484
transform 1 0 48944 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1666464484
transform 1 0 54924 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1666464484
transform 1 0 4048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1666464484
transform 1 0 10028 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1666464484
transform 1 0 16008 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1666464484
transform 1 0 21988 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1666464484
transform 1 0 27968 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1666464484
transform 1 0 33948 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1666464484
transform 1 0 39928 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1666464484
transform 1 0 45908 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1666464484
transform 1 0 51888 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1666464484
transform 1 0 57868 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1666464484
transform 1 0 7084 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1666464484
transform 1 0 13064 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1666464484
transform 1 0 19044 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1666464484
transform 1 0 25024 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1666464484
transform 1 0 31004 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1666464484
transform 1 0 36984 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1666464484
transform 1 0 42964 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1666464484
transform 1 0 48944 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1666464484
transform 1 0 54924 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1666464484
transform 1 0 4048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1666464484
transform 1 0 10028 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1666464484
transform 1 0 16008 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1666464484
transform 1 0 21988 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1666464484
transform 1 0 27968 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1666464484
transform 1 0 33948 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1666464484
transform 1 0 39928 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1666464484
transform 1 0 45908 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1666464484
transform 1 0 51888 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1666464484
transform 1 0 57868 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1666464484
transform 1 0 4048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1666464484
transform 1 0 6992 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1666464484
transform 1 0 9936 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1666464484
transform 1 0 12880 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1666464484
transform 1 0 15824 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1666464484
transform 1 0 18768 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1666464484
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1666464484
transform 1 0 24656 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1666464484
transform 1 0 27600 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1666464484
transform 1 0 30544 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1666464484
transform 1 0 33488 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1666464484
transform 1 0 36432 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1666464484
transform 1 0 39376 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1666464484
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1666464484
transform 1 0 45264 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1666464484
transform 1 0 48208 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1666464484
transform 1 0 51152 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1666464484
transform 1 0 54096 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1666464484
transform 1 0 57040 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _157_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26864 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _158_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23920 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _159_
timestamp 1666464484
transform 1 0 30268 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1666464484
transform 1 0 37352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1666464484
transform -1 0 36800 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1666464484
transform 1 0 34224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1666464484
transform -1 0 36984 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1666464484
transform 1 0 37260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1666464484
transform -1 0 35236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1666464484
transform 1 0 32936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1666464484
transform -1 0 36800 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1666464484
transform 1 0 30544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _170_
timestamp 1666464484
transform 1 0 29992 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1666464484
transform 1 0 30820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1666464484
transform 1 0 30728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1666464484
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1666464484
transform 1 0 28980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1666464484
transform 1 0 29992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1666464484
transform -1 0 29624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1666464484
transform 1 0 28244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1666464484
transform 1 0 25944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1666464484
transform 1 0 24196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1666464484
transform -1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _181_
timestamp 1666464484
transform 1 0 26680 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1666464484
transform 1 0 23920 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1666464484
transform 1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1666464484
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1666464484
transform 1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1666464484
transform 1 0 27600 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1666464484
transform -1 0 27048 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1666464484
transform -1 0 22264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1666464484
transform 1 0 22264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1666464484
transform 1 0 22908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1666464484
transform 1 0 23920 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1666464484
transform 1 0 24564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _193_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 36432 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _194_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34960 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _195_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 35328 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _196_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29992 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _197_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 36248 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _198_
timestamp 1666464484
transform -1 0 35328 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _199_
timestamp 1666464484
transform -1 0 30268 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _200_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34776 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _201_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34316 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _202_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32844 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _203_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31740 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _204_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 33764 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _205_
timestamp 1666464484
transform 1 0 31924 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _206_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29900 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _207_
timestamp 1666464484
transform -1 0 29808 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _208_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29072 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _209_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34592 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _210_
timestamp 1666464484
transform 1 0 28336 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _211_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28428 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _212_
timestamp 1666464484
transform -1 0 28428 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _213_
timestamp 1666464484
transform -1 0 45724 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _214_
timestamp 1666464484
transform 1 0 44620 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _215_
timestamp 1666464484
transform -1 0 44896 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _216_
timestamp 1666464484
transform -1 0 40664 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _217_
timestamp 1666464484
transform 1 0 44528 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _218_
timestamp 1666464484
transform -1 0 44160 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _219_
timestamp 1666464484
transform -1 0 39560 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _220_
timestamp 1666464484
transform -1 0 43792 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _221_
timestamp 1666464484
transform -1 0 43148 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _222_
timestamp 1666464484
transform 1 0 41952 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _223_
timestamp 1666464484
transform 1 0 40664 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _224_
timestamp 1666464484
transform -1 0 42320 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _225_
timestamp 1666464484
transform 1 0 40756 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _226_
timestamp 1666464484
transform -1 0 39008 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _227_
timestamp 1666464484
transform -1 0 39468 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _228_
timestamp 1666464484
transform 1 0 38088 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _229_
timestamp 1666464484
transform -1 0 44252 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _230_
timestamp 1666464484
transform 1 0 37352 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _231_
timestamp 1666464484
transform 1 0 37720 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _232_
timestamp 1666464484
transform -1 0 35788 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _233_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34868 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _234_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27876 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _235_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1666464484
transform -1 0 33764 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _237_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31740 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _238_
timestamp 1666464484
transform 1 0 31464 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _239_
timestamp 1666464484
transform 1 0 30728 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1666464484
transform -1 0 39192 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _241_
timestamp 1666464484
transform 1 0 41124 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _242_
timestamp 1666464484
transform 1 0 40204 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _243_
timestamp 1666464484
transform 1 0 40020 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _244_
timestamp 1666464484
transform 1 0 23644 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _245_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23828 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _246_
timestamp 1666464484
transform -1 0 24288 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1666464484
transform -1 0 23552 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _248_
timestamp 1666464484
transform -1 0 24104 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _249_
timestamp 1666464484
transform -1 0 32936 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _250_
timestamp 1666464484
transform 1 0 32200 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _251_
timestamp 1666464484
transform 1 0 34132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _252_
timestamp 1666464484
transform 1 0 33120 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _253_
timestamp 1666464484
transform 1 0 32844 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _254_
timestamp 1666464484
transform -1 0 42136 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _255_
timestamp 1666464484
transform 1 0 40940 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _256_
timestamp 1666464484
transform 1 0 42320 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _257_
timestamp 1666464484
transform 1 0 41952 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _258_
timestamp 1666464484
transform 1 0 41032 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _259_
timestamp 1666464484
transform 1 0 25300 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1666464484
transform 1 0 25484 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _261_
timestamp 1666464484
transform -1 0 25668 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1666464484
transform -1 0 24840 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _263_
timestamp 1666464484
transform 1 0 25024 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _264_
timestamp 1666464484
transform 1 0 31924 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _265_
timestamp 1666464484
transform 1 0 32660 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _266_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30176 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _267_
timestamp 1666464484
transform 1 0 30360 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _268_
timestamp 1666464484
transform -1 0 31096 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _269_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31556 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _270_
timestamp 1666464484
transform -1 0 43792 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _271_
timestamp 1666464484
transform -1 0 42136 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _272_
timestamp 1666464484
transform 1 0 39008 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _273_
timestamp 1666464484
transform 1 0 41032 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _274_
timestamp 1666464484
transform -1 0 40204 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _275_
timestamp 1666464484
transform 1 0 39836 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _276_
timestamp 1666464484
transform -1 0 26680 0 1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1666464484
transform 1 0 26220 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _278_
timestamp 1666464484
transform -1 0 27140 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _279_
timestamp 1666464484
transform -1 0 26312 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _280_
timestamp 1666464484
transform -1 0 26956 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _281_
timestamp 1666464484
transform -1 0 28704 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _282_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29072 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _283_
timestamp 1666464484
transform 1 0 28336 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _284_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27416 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _285_
timestamp 1666464484
transform 1 0 32844 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _286_
timestamp 1666464484
transform 1 0 33764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _287_
timestamp 1666464484
transform -1 0 27600 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _288_
timestamp 1666464484
transform 1 0 38088 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _289_
timestamp 1666464484
transform -1 0 38180 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _290_
timestamp 1666464484
transform 1 0 36340 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _291_
timestamp 1666464484
transform 1 0 42780 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _292_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 43700 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _293_
timestamp 1666464484
transform 1 0 36248 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _294_
timestamp 1666464484
transform 1 0 35972 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _295_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29900 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _296_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28888 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _519__194 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 25576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25300 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _520__195
timestamp 1666464484
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _520_
timestamp 1666464484
transform 1 0 25852 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _521__196
timestamp 1666464484
transform 1 0 23276 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _521_
timestamp 1666464484
transform 1 0 25852 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _522_
timestamp 1666464484
transform 1 0 23552 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _522__197
timestamp 1666464484
transform 1 0 22264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _523_
timestamp 1666464484
transform 1 0 25484 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _523__198
timestamp 1666464484
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _524_
timestamp 1666464484
transform 1 0 25852 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _524__199
timestamp 1666464484
transform 1 0 25208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _525_
timestamp 1666464484
transform 1 0 27692 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _525__200
timestamp 1666464484
transform 1 0 26036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _526__201
timestamp 1666464484
transform 1 0 27508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _526_
timestamp 1666464484
transform 1 0 27600 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _527__202
timestamp 1666464484
transform 1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _527_
timestamp 1666464484
transform 1 0 28244 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _528__203
timestamp 1666464484
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _528_
timestamp 1666464484
transform 1 0 27876 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _529_
timestamp 1666464484
transform 1 0 26588 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _529__204
timestamp 1666464484
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _530_
timestamp 1666464484
transform 1 0 25576 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _530__205
timestamp 1666464484
transform 1 0 23552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _531_
timestamp 1666464484
transform 1 0 28428 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _531__206
timestamp 1666464484
transform 1 0 23920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _532__207
timestamp 1666464484
transform 1 0 28336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _532_
timestamp 1666464484
transform 1 0 28888 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _533__208
timestamp 1666464484
transform 1 0 28704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _533_
timestamp 1666464484
transform 1 0 28888 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _534__209
timestamp 1666464484
transform -1 0 29716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _534_
timestamp 1666464484
transform 1 0 28704 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _535__210
timestamp 1666464484
transform -1 0 30360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _535_
timestamp 1666464484
transform 1 0 29992 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _536__211
timestamp 1666464484
transform 1 0 29624 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _536_
timestamp 1666464484
transform 1 0 30268 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _537__212
timestamp 1666464484
transform -1 0 36432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _537_
timestamp 1666464484
transform -1 0 32752 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _538_
timestamp 1666464484
transform 1 0 31280 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _538__213
timestamp 1666464484
transform -1 0 31556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _539__214
timestamp 1666464484
transform -1 0 31556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _539_
timestamp 1666464484
transform 1 0 31004 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _540__215
timestamp 1666464484
transform -1 0 32200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _540_
timestamp 1666464484
transform 1 0 31464 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _541__216
timestamp 1666464484
transform -1 0 35880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _541_
timestamp 1666464484
transform -1 0 33488 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _542__217
timestamp 1666464484
transform 1 0 32292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _542_
timestamp 1666464484
transform -1 0 33764 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _543_
timestamp 1666464484
transform 1 0 33580 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _543__218
timestamp 1666464484
transform 1 0 32568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _544__219
timestamp 1666464484
transform 1 0 33212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _544_
timestamp 1666464484
transform -1 0 34592 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _545__220
timestamp 1666464484
transform -1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _545_
timestamp 1666464484
transform -1 0 35788 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _546__221
timestamp 1666464484
transform -1 0 37444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _546_
timestamp 1666464484
transform -1 0 35696 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _547__222
timestamp 1666464484
transform 1 0 34132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _547_
timestamp 1666464484
transform 1 0 34224 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _548__223
timestamp 1666464484
transform 1 0 35880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _548_
timestamp 1666464484
transform -1 0 36156 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _549__224
timestamp 1666464484
transform -1 0 37536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _549_
timestamp 1666464484
transform -1 0 36156 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _550_
timestamp 1666464484
transform 1 0 34040 0 -1 52224
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _550__225
timestamp 1666464484
transform -1 0 34500 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4324 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform -1 0 27784 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform -1 0 29716 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 32752 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1666464484
transform 1 0 35420 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1666464484
transform -1 0 35052 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1666464484
transform 1 0 36708 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1666464484
transform 1 0 37996 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1666464484
transform 1 0 38732 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1666464484
transform -1 0 40388 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1666464484
transform 1 0 44988 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1666464484
transform 1 0 42872 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1666464484
transform 1 0 46828 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1666464484
transform -1 0 46000 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1666464484
transform 1 0 47012 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1666464484
transform 1 0 48484 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1666464484
transform 1 0 49772 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 51428 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 52532 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1666464484
transform 1 0 54372 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1666464484
transform -1 0 55660 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  macro_15_37
timestamp 1666464484
transform -1 0 50968 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_38
timestamp 1666464484
transform -1 0 52440 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_39
timestamp 1666464484
transform -1 0 53728 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_40
timestamp 1666464484
transform -1 0 54648 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_41
timestamp 1666464484
transform -1 0 56304 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_42
timestamp 1666464484
transform -1 0 6808 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_43
timestamp 1666464484
transform -1 0 8188 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_44
timestamp 1666464484
transform -1 0 9568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_45
timestamp 1666464484
transform -1 0 30268 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_46
timestamp 1666464484
transform 1 0 30084 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_47
timestamp 1666464484
transform -1 0 34500 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_48
timestamp 1666464484
transform -1 0 35420 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_49
timestamp 1666464484
transform -1 0 37536 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_50
timestamp 1666464484
transform -1 0 41308 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_51
timestamp 1666464484
transform -1 0 38548 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_52
timestamp 1666464484
transform -1 0 45080 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_53
timestamp 1666464484
transform -1 0 41952 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_54
timestamp 1666464484
transform -1 0 43516 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_55
timestamp 1666464484
transform -1 0 46460 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_56
timestamp 1666464484
transform -1 0 47012 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_57
timestamp 1666464484
transform -1 0 47656 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_58
timestamp 1666464484
transform -1 0 49036 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_59
timestamp 1666464484
transform -1 0 50324 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_60
timestamp 1666464484
transform -1 0 51612 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_61
timestamp 1666464484
transform -1 0 53084 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_62
timestamp 1666464484
transform -1 0 53728 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_63
timestamp 1666464484
transform -1 0 55292 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_64
timestamp 1666464484
transform -1 0 56488 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_65
timestamp 1666464484
transform -1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_66
timestamp 1666464484
transform 1 0 16376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_67
timestamp 1666464484
transform 1 0 17296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_68
timestamp 1666464484
transform -1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_69
timestamp 1666464484
transform 1 0 17020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_70
timestamp 1666464484
transform 1 0 17940 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_71
timestamp 1666464484
transform -1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_72
timestamp 1666464484
transform 1 0 17664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_73
timestamp 1666464484
transform 1 0 18584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_74
timestamp 1666464484
transform -1 0 20148 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_75
timestamp 1666464484
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_76
timestamp 1666464484
transform 1 0 19596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_77
timestamp 1666464484
transform -1 0 20976 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_78
timestamp 1666464484
transform 1 0 20240 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_79
timestamp 1666464484
transform 1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_80
timestamp 1666464484
transform -1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_81
timestamp 1666464484
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_82
timestamp 1666464484
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_83
timestamp 1666464484
transform 1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_84
timestamp 1666464484
transform -1 0 22908 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_85
timestamp 1666464484
transform 1 0 19320 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_86
timestamp 1666464484
transform -1 0 23460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_87
timestamp 1666464484
transform 1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_88
timestamp 1666464484
transform 1 0 21988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_89
timestamp 1666464484
transform 1 0 23276 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_90
timestamp 1666464484
transform 1 0 21528 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_91
timestamp 1666464484
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_92
timestamp 1666464484
transform 1 0 23920 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_93
timestamp 1666464484
transform 1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_94
timestamp 1666464484
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_95
timestamp 1666464484
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_96
timestamp 1666464484
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_97
timestamp 1666464484
transform -1 0 38272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_98
timestamp 1666464484
transform -1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_99
timestamp 1666464484
transform -1 0 38916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_100
timestamp 1666464484
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_101
timestamp 1666464484
transform -1 0 38088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_102
timestamp 1666464484
transform -1 0 39928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_103
timestamp 1666464484
transform -1 0 38732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_104
timestamp 1666464484
transform -1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_105
timestamp 1666464484
transform -1 0 38180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_106
timestamp 1666464484
transform -1 0 39376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_107
timestamp 1666464484
transform -1 0 40572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_108
timestamp 1666464484
transform -1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_109
timestamp 1666464484
transform -1 0 41216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_110
timestamp 1666464484
transform -1 0 38916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_111
timestamp 1666464484
transform -1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_112
timestamp 1666464484
transform -1 0 41860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_113
timestamp 1666464484
transform -1 0 40480 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_114
timestamp 1666464484
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_115
timestamp 1666464484
transform -1 0 41124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_116
timestamp 1666464484
transform -1 0 42044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_117
timestamp 1666464484
transform -1 0 42872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_118
timestamp 1666464484
transform -1 0 41768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_119
timestamp 1666464484
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_120
timestamp 1666464484
transform -1 0 42412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_121
timestamp 1666464484
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_122
timestamp 1666464484
transform -1 0 43516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_123
timestamp 1666464484
transform -1 0 44160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_124
timestamp 1666464484
transform -1 0 43056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_125
timestamp 1666464484
transform -1 0 44804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_126
timestamp 1666464484
transform -1 0 44160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_127
timestamp 1666464484
transform -1 0 43700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_128
timestamp 1666464484
transform -1 0 44804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_129
timestamp 1666464484
transform -1 0 45816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_130
timestamp 1666464484
transform -1 0 44436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_131
timestamp 1666464484
transform -1 0 45448 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_132
timestamp 1666464484
transform -1 0 46460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_133
timestamp 1666464484
transform -1 0 46092 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_134
timestamp 1666464484
transform -1 0 47104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_135
timestamp 1666464484
transform -1 0 46736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_136
timestamp 1666464484
transform -1 0 47748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_137
timestamp 1666464484
transform -1 0 46460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_138
timestamp 1666464484
transform -1 0 47380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_139
timestamp 1666464484
transform -1 0 47104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_140
timestamp 1666464484
transform -1 0 48024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_141
timestamp 1666464484
transform -1 0 48760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_142
timestamp 1666464484
transform -1 0 49404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_143
timestamp 1666464484
transform -1 0 48668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_144
timestamp 1666464484
transform -1 0 50048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_145
timestamp 1666464484
transform -1 0 48576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_146
timestamp 1666464484
transform -1 0 49496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_147
timestamp 1666464484
transform -1 0 50692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_148
timestamp 1666464484
transform -1 0 50140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_149
timestamp 1666464484
transform -1 0 49680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_150
timestamp 1666464484
transform -1 0 50784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_151
timestamp 1666464484
transform -1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_152
timestamp 1666464484
transform -1 0 50508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_153
timestamp 1666464484
transform -1 0 51428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_154
timestamp 1666464484
transform -1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_155
timestamp 1666464484
transform -1 0 52072 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_156
timestamp 1666464484
transform -1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_157
timestamp 1666464484
transform -1 0 52716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_158
timestamp 1666464484
transform -1 0 53636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_159
timestamp 1666464484
transform -1 0 52440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_160
timestamp 1666464484
transform -1 0 53360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_161
timestamp 1666464484
transform -1 0 8004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_162
timestamp 1666464484
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_163
timestamp 1666464484
transform -1 0 8924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_164
timestamp 1666464484
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_165
timestamp 1666464484
transform -1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_166
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_167
timestamp 1666464484
transform 1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_168
timestamp 1666464484
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_169
timestamp 1666464484
transform 1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_170
timestamp 1666464484
transform -1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_171
timestamp 1666464484
transform 1 0 10672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_172
timestamp 1666464484
transform 1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_173
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_174
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_175
timestamp 1666464484
transform 1 0 11960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_176
timestamp 1666464484
transform -1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_177
timestamp 1666464484
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_178
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_179
timestamp 1666464484
transform 1 0 12420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_180
timestamp 1666464484
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_181
timestamp 1666464484
transform 1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_182
timestamp 1666464484
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_183
timestamp 1666464484
transform 1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_184
timestamp 1666464484
transform -1 0 14996 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_185
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_186
timestamp 1666464484
transform 1 0 14720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_187
timestamp 1666464484
transform -1 0 15824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_188
timestamp 1666464484
transform 1 0 14720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_189
timestamp 1666464484
transform 1 0 15364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_190
timestamp 1666464484
transform 1 0 15364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_191
timestamp 1666464484
transform -1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_192
timestamp 1666464484
transform 1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_193
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_226
timestamp 1666464484
transform -1 0 4968 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_227
timestamp 1666464484
transform -1 0 6164 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_228
timestamp 1666464484
transform -1 0 7544 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_229
timestamp 1666464484
transform -1 0 8924 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_230
timestamp 1666464484
transform -1 0 10580 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_231
timestamp 1666464484
transform -1 0 11684 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_232
timestamp 1666464484
transform -1 0 13248 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_233
timestamp 1666464484
transform -1 0 14444 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_234
timestamp 1666464484
transform -1 0 16560 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_235
timestamp 1666464484
transform -1 0 17204 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_236
timestamp 1666464484
transform -1 0 18584 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_237
timestamp 1666464484
transform -1 0 20148 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_238
timestamp 1666464484
transform -1 0 21528 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_239
timestamp 1666464484
transform -1 0 22908 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_240
timestamp 1666464484
transform 1 0 21252 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_241
timestamp 1666464484
transform 1 0 22724 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_242
timestamp 1666464484
transform -1 0 27048 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_243
timestamp 1666464484
transform 1 0 27508 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_244
timestamp 1666464484
transform -1 0 30360 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_245
timestamp 1666464484
transform -1 0 31188 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_246
timestamp 1666464484
transform -1 0 32660 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_247
timestamp 1666464484
transform -1 0 35972 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_248
timestamp 1666464484
transform -1 0 36064 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_249
timestamp 1666464484
transform -1 0 36708 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_250
timestamp 1666464484
transform -1 0 38088 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_251
timestamp 1666464484
transform -1 0 44436 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_252
timestamp 1666464484
transform -1 0 43516 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_253
timestamp 1666464484
transform -1 0 42780 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_254
timestamp 1666464484
transform -1 0 46644 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_255
timestamp 1666464484
transform -1 0 46368 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_256
timestamp 1666464484
transform -1 0 47748 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_257
timestamp 1666464484
transform -1 0 48392 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_15_258
timestamp 1666464484
transform -1 0 49680 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1666464484
transform -1 0 5520 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1666464484
transform -1 0 19412 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1666464484
transform -1 0 20700 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1666464484
transform -1 0 22356 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1666464484
transform -1 0 23460 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1666464484
transform 1 0 24932 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1666464484
transform 1 0 25852 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1666464484
transform 1 0 27876 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1666464484
transform -1 0 28980 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1666464484
transform -1 0 11040 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1666464484
transform -1 0 12420 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1666464484
transform -1 0 13800 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1666464484
transform -1 0 15180 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1666464484
transform -1 0 16560 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1666464484
transform -1 0 17940 0 -1 57664
box -38 -48 406 592
<< labels >>
flabel metal2 s 3698 59200 3754 60000 0 FreeSans 224 90 0 0 io_active
port 0 nsew signal input
flabel metal2 s 4158 59200 4214 60000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 17958 59200 18014 60000 0 FreeSans 224 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s 19338 59200 19394 60000 0 FreeSans 224 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal2 s 20718 59200 20774 60000 0 FreeSans 224 90 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 22098 59200 22154 60000 0 FreeSans 224 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 23478 59200 23534 60000 0 FreeSans 224 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal2 s 24858 59200 24914 60000 0 FreeSans 224 90 0 0 io_in[15]
port 7 nsew signal input
flabel metal2 s 26238 59200 26294 60000 0 FreeSans 224 90 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 27618 59200 27674 60000 0 FreeSans 224 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 28998 59200 29054 60000 0 FreeSans 224 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 30378 59200 30434 60000 0 FreeSans 224 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal2 s 5538 59200 5594 60000 0 FreeSans 224 90 0 0 io_in[1]
port 12 nsew signal input
flabel metal2 s 31758 59200 31814 60000 0 FreeSans 224 90 0 0 io_in[20]
port 13 nsew signal input
flabel metal2 s 33138 59200 33194 60000 0 FreeSans 224 90 0 0 io_in[21]
port 14 nsew signal input
flabel metal2 s 34518 59200 34574 60000 0 FreeSans 224 90 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 35898 59200 35954 60000 0 FreeSans 224 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 37278 59200 37334 60000 0 FreeSans 224 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 38658 59200 38714 60000 0 FreeSans 224 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 40038 59200 40094 60000 0 FreeSans 224 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal2 s 41418 59200 41474 60000 0 FreeSans 224 90 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 42798 59200 42854 60000 0 FreeSans 224 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 44178 59200 44234 60000 0 FreeSans 224 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 6918 59200 6974 60000 0 FreeSans 224 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal2 s 45558 59200 45614 60000 0 FreeSans 224 90 0 0 io_in[30]
port 24 nsew signal input
flabel metal2 s 46938 59200 46994 60000 0 FreeSans 224 90 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 48318 59200 48374 60000 0 FreeSans 224 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal2 s 49698 59200 49754 60000 0 FreeSans 224 90 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 51078 59200 51134 60000 0 FreeSans 224 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 52458 59200 52514 60000 0 FreeSans 224 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal2 s 53838 59200 53894 60000 0 FreeSans 224 90 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 55218 59200 55274 60000 0 FreeSans 224 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 8298 59200 8354 60000 0 FreeSans 224 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal2 s 9678 59200 9734 60000 0 FreeSans 224 90 0 0 io_in[4]
port 33 nsew signal input
flabel metal2 s 11058 59200 11114 60000 0 FreeSans 224 90 0 0 io_in[5]
port 34 nsew signal input
flabel metal2 s 12438 59200 12494 60000 0 FreeSans 224 90 0 0 io_in[6]
port 35 nsew signal input
flabel metal2 s 13818 59200 13874 60000 0 FreeSans 224 90 0 0 io_in[7]
port 36 nsew signal input
flabel metal2 s 15198 59200 15254 60000 0 FreeSans 224 90 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 16578 59200 16634 60000 0 FreeSans 224 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 4618 59200 4674 60000 0 FreeSans 224 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal2 s 18418 59200 18474 60000 0 FreeSans 224 90 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal2 s 19798 59200 19854 60000 0 FreeSans 224 90 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal2 s 21178 59200 21234 60000 0 FreeSans 224 90 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal2 s 22558 59200 22614 60000 0 FreeSans 224 90 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal2 s 23938 59200 23994 60000 0 FreeSans 224 90 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 25318 59200 25374 60000 0 FreeSans 224 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal2 s 26698 59200 26754 60000 0 FreeSans 224 90 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 28078 59200 28134 60000 0 FreeSans 224 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 29458 59200 29514 60000 0 FreeSans 224 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 30838 59200 30894 60000 0 FreeSans 224 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal2 s 5998 59200 6054 60000 0 FreeSans 224 90 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal2 s 32218 59200 32274 60000 0 FreeSans 224 90 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal2 s 33598 59200 33654 60000 0 FreeSans 224 90 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 34978 59200 35034 60000 0 FreeSans 224 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 36358 59200 36414 60000 0 FreeSans 224 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 37738 59200 37794 60000 0 FreeSans 224 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal2 s 39118 59200 39174 60000 0 FreeSans 224 90 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal2 s 40498 59200 40554 60000 0 FreeSans 224 90 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 41878 59200 41934 60000 0 FreeSans 224 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal2 s 43258 59200 43314 60000 0 FreeSans 224 90 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal2 s 44638 59200 44694 60000 0 FreeSans 224 90 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 7378 59200 7434 60000 0 FreeSans 224 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal2 s 46018 59200 46074 60000 0 FreeSans 224 90 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal2 s 47398 59200 47454 60000 0 FreeSans 224 90 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal2 s 48778 59200 48834 60000 0 FreeSans 224 90 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal2 s 50158 59200 50214 60000 0 FreeSans 224 90 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal2 s 51538 59200 51594 60000 0 FreeSans 224 90 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal2 s 52918 59200 52974 60000 0 FreeSans 224 90 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal2 s 54298 59200 54354 60000 0 FreeSans 224 90 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal2 s 55678 59200 55734 60000 0 FreeSans 224 90 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 8758 59200 8814 60000 0 FreeSans 224 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal2 s 10138 59200 10194 60000 0 FreeSans 224 90 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal2 s 11518 59200 11574 60000 0 FreeSans 224 90 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal2 s 12898 59200 12954 60000 0 FreeSans 224 90 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 14278 59200 14334 60000 0 FreeSans 224 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 15658 59200 15714 60000 0 FreeSans 224 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 17038 59200 17094 60000 0 FreeSans 224 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal2 s 5078 59200 5134 60000 0 FreeSans 224 90 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal2 s 18878 59200 18934 60000 0 FreeSans 224 90 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal2 s 20258 59200 20314 60000 0 FreeSans 224 90 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal2 s 21638 59200 21694 60000 0 FreeSans 224 90 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal2 s 23018 59200 23074 60000 0 FreeSans 224 90 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal2 s 24398 59200 24454 60000 0 FreeSans 224 90 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal2 s 25778 59200 25834 60000 0 FreeSans 224 90 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal2 s 27158 59200 27214 60000 0 FreeSans 224 90 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 28538 59200 28594 60000 0 FreeSans 224 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal2 s 29918 59200 29974 60000 0 FreeSans 224 90 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal2 s 31298 59200 31354 60000 0 FreeSans 224 90 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 6458 59200 6514 60000 0 FreeSans 224 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 32678 59200 32734 60000 0 FreeSans 224 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal2 s 34058 59200 34114 60000 0 FreeSans 224 90 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 35438 59200 35494 60000 0 FreeSans 224 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal2 s 36818 59200 36874 60000 0 FreeSans 224 90 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 38198 59200 38254 60000 0 FreeSans 224 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 39578 59200 39634 60000 0 FreeSans 224 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal2 s 40958 59200 41014 60000 0 FreeSans 224 90 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 42338 59200 42394 60000 0 FreeSans 224 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 43718 59200 43774 60000 0 FreeSans 224 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal2 s 45098 59200 45154 60000 0 FreeSans 224 90 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 7838 59200 7894 60000 0 FreeSans 224 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal2 s 46478 59200 46534 60000 0 FreeSans 224 90 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal2 s 47858 59200 47914 60000 0 FreeSans 224 90 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal2 s 49238 59200 49294 60000 0 FreeSans 224 90 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal2 s 50618 59200 50674 60000 0 FreeSans 224 90 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal2 s 51998 59200 52054 60000 0 FreeSans 224 90 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal2 s 53378 59200 53434 60000 0 FreeSans 224 90 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 54758 59200 54814 60000 0 FreeSans 224 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal2 s 56138 59200 56194 60000 0 FreeSans 224 90 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal2 s 9218 59200 9274 60000 0 FreeSans 224 90 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal2 s 10598 59200 10654 60000 0 FreeSans 224 90 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 11978 59200 12034 60000 0 FreeSans 224 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 13358 59200 13414 60000 0 FreeSans 224 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal2 s 14738 59200 14794 60000 0 FreeSans 224 90 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 16118 59200 16174 60000 0 FreeSans 224 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal2 s 17498 59200 17554 60000 0 FreeSans 224 90 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 115 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 116 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 117 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 118 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 119 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 120 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 121 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 122 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 123 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 124 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 125 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 126 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 127 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 128 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 129 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 130 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 131 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 132 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 133 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 134 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 135 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 136 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 137 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 138 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 139 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 140 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 141 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 142 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 143 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 144 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 145 nsew signal input
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 146 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 147 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 148 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 149 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 150 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 151 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 152 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 153 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 154 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 155 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 156 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 157 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 158 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 159 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 160 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 161 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 162 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 163 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 164 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 165 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 166 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 167 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 168 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 169 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 170 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 171 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 172 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 173 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 174 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 175 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 176 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 177 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 178 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 179 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 180 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 181 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 182 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 183 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 184 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 185 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 186 nsew signal input
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 187 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 188 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 189 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 190 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 191 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 192 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 193 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 194 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 195 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 196 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 197 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 198 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 199 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 200 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 201 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 202 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 203 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 204 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 205 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 206 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 207 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 208 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 209 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 210 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 211 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 212 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 213 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 214 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 215 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 216 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 217 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 218 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 219 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 220 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 221 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 222 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 223 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 224 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 225 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 226 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 227 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 228 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 229 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 230 nsew signal input
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 231 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 232 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 233 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 234 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 235 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 236 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 237 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 238 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 239 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 240 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 241 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 242 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 243 nsew signal tristate
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 244 nsew signal tristate
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 245 nsew signal tristate
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 246 nsew signal tristate
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 247 nsew signal tristate
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 248 nsew signal tristate
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 249 nsew signal tristate
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 250 nsew signal tristate
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 251 nsew signal tristate
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 252 nsew signal tristate
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 253 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 254 nsew signal tristate
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 255 nsew signal tristate
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 256 nsew signal tristate
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 257 nsew signal tristate
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 258 nsew signal tristate
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 259 nsew signal tristate
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 260 nsew signal tristate
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 261 nsew signal tristate
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 262 nsew signal tristate
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 263 nsew signal tristate
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 264 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 265 nsew signal tristate
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 266 nsew signal tristate
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 267 nsew signal tristate
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 268 nsew signal tristate
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 269 nsew signal tristate
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 270 nsew signal tristate
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 271 nsew signal tristate
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 272 nsew signal tristate
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 273 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 274 nsew signal tristate
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 275 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 276 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 277 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 278 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 279 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 280 nsew signal tristate
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 281 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 282 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 283 nsew signal tristate
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 284 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 285 nsew signal tristate
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 286 nsew signal tristate
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 287 nsew signal tristate
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 288 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 289 nsew signal tristate
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 290 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 291 nsew signal tristate
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 292 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 293 nsew signal tristate
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 294 nsew signal tristate
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 295 nsew signal tristate
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 296 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 297 nsew signal tristate
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 298 nsew signal tristate
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 299 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 300 nsew signal tristate
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 301 nsew signal tristate
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 302 nsew signal tristate
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 303 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 304 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 305 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 306 nsew signal tristate
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 307 nsew signal tristate
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 308 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 309 nsew signal tristate
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 310 nsew signal tristate
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 311 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 312 nsew signal tristate
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 313 nsew signal tristate
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 314 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 315 nsew signal tristate
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 316 nsew signal tristate
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 317 nsew signal tristate
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 318 nsew signal tristate
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 319 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 320 nsew signal tristate
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 321 nsew signal tristate
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 322 nsew signal tristate
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 323 nsew signal tristate
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 324 nsew signal tristate
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 325 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 326 nsew signal tristate
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 327 nsew signal tristate
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 328 nsew signal tristate
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 329 nsew signal tristate
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 330 nsew signal tristate
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 331 nsew signal tristate
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 332 nsew signal tristate
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 333 nsew signal tristate
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 334 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 335 nsew signal tristate
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 336 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 337 nsew signal tristate
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 338 nsew signal tristate
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 339 nsew signal tristate
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 340 nsew signal tristate
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 341 nsew signal tristate
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 342 nsew signal tristate
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 343 nsew signal tristate
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 344 nsew signal tristate
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 345 nsew signal tristate
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 346 nsew signal tristate
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 347 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 348 nsew signal tristate
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 349 nsew signal tristate
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 350 nsew signal tristate
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 351 nsew signal tristate
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 352 nsew signal tristate
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 353 nsew signal tristate
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 354 nsew signal tristate
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 355 nsew signal tristate
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 356 nsew signal tristate
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 357 nsew signal tristate
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 358 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 359 nsew signal tristate
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 360 nsew signal tristate
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 361 nsew signal tristate
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 362 nsew signal tristate
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 363 nsew signal tristate
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 364 nsew signal tristate
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 365 nsew signal tristate
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 366 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 367 nsew signal tristate
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 368 nsew signal tristate
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 369 nsew signal tristate
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 370 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 371 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 372 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 373 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 374 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 375 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 376 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 377 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 378 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 379 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 380 nsew signal input
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 381 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 382 nsew signal input
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 383 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 384 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 385 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 386 nsew signal input
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 387 nsew signal input
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 388 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 389 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 390 nsew signal input
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 391 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 392 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 393 nsew signal input
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 394 nsew signal input
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 395 nsew signal input
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 396 nsew signal input
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 397 nsew signal input
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 398 nsew signal input
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 399 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 400 nsew signal input
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 401 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 402 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 403 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 404 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 405 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 406 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 407 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 408 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 409 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 410 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 411 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 412 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 413 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 414 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 415 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 416 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 417 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 418 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 419 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 420 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 421 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 422 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 423 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 424 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 425 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 426 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 427 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 428 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 429 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 430 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 431 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 432 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 433 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 434 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 435 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 436 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 437 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 438 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 439 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 440 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 441 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 442 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 443 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 444 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 445 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 446 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 447 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 448 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 449 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 450 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 451 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 452 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 453 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 454 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 455 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 456 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 457 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 458 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 459 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 460 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 461 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 462 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 463 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 464 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 465 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 466 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 467 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 468 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 469 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 470 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 471 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 472 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 473 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 474 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 475 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 476 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 477 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 478 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 479 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 480 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 481 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 482 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 483 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 484 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 485 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 486 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 487 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 488 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 489 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 490 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 491 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 492 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 493 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 494 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 495 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 496 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 497 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 498 nsew signal input
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 500 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 500 nsew ground bidirectional
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wb_clk_i
port 501 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wb_rst_i
port 502 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 503 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 504 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 505 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 506 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 507 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 508 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 509 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 510 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 511 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 512 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 513 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 514 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 515 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 516 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 517 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 518 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 519 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 520 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 521 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 522 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 523 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 524 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 525 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 526 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 527 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 528 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 529 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 530 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 531 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 532 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 533 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 534 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 535 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 536 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 537 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 538 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 539 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 540 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 541 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 542 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 543 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 544 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 545 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 546 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 547 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 548 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 549 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 550 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 551 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 552 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 553 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 554 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 555 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 556 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 557 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 558 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 559 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 560 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 561 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 562 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 563 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 564 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 565 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 566 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 567 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 568 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 569 nsew signal tristate
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 570 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 571 nsew signal tristate
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 572 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 573 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 574 nsew signal tristate
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 575 nsew signal tristate
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 576 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 577 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 578 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 579 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 580 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 581 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 582 nsew signal tristate
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 583 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 584 nsew signal tristate
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 585 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 586 nsew signal tristate
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 587 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 588 nsew signal tristate
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 589 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 590 nsew signal tristate
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 591 nsew signal tristate
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 592 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 593 nsew signal tristate
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 594 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 595 nsew signal tristate
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 596 nsew signal tristate
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 597 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 598 nsew signal tristate
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 599 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 600 nsew signal tristate
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 601 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 602 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 603 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 604 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 605 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_we_i
port 606 nsew signal input
rlabel metal1 29992 57120 29992 57120 0 vccd1
rlabel metal1 29992 57664 29992 57664 0 vssd1
rlabel metal2 34454 54400 34454 54400 0 _000_
rlabel metal2 35006 55590 35006 55590 0 _001_
rlabel metal1 34730 55828 34730 55828 0 _002_
rlabel metal1 28658 55794 28658 55794 0 _003_
rlabel metal1 35190 54060 35190 54060 0 _004_
rlabel metal1 30498 54060 30498 54060 0 _005_
rlabel metal2 29026 54128 29026 54128 0 _006_
rlabel metal1 33764 54502 33764 54502 0 _007_
rlabel metal1 33488 54298 33488 54298 0 _008_
rlabel metal1 32614 54502 32614 54502 0 _009_
rlabel metal2 32430 54842 32430 54842 0 _010_
rlabel metal2 32614 54162 32614 54162 0 _011_
rlabel metal1 31372 54638 31372 54638 0 _012_
rlabel metal1 29256 55318 29256 55318 0 _013_
rlabel metal1 29302 54298 29302 54298 0 _014_
rlabel via1 28658 55709 28658 55709 0 _015_
rlabel metal1 33806 55386 33806 55386 0 _016_
rlabel metal1 27968 56338 27968 56338 0 _017_
rlabel metal2 28474 55522 28474 55522 0 _018_
rlabel metal1 27876 56474 27876 56474 0 _019_
rlabel metal1 45310 55726 45310 55726 0 _020_
rlabel metal1 44620 55930 44620 55930 0 _021_
rlabel via1 40618 55675 40618 55675 0 _022_
rlabel metal1 38088 56202 38088 56202 0 _023_
rlabel metal1 44298 54706 44298 54706 0 _024_
rlabel metal1 39330 54740 39330 54740 0 _025_
rlabel metal1 38824 55386 38824 55386 0 _026_
rlabel metal1 42826 54230 42826 54230 0 _027_
rlabel metal2 42458 54332 42458 54332 0 _028_
rlabel metal2 41998 54774 41998 54774 0 _029_
rlabel metal2 41262 54842 41262 54842 0 _030_
rlabel metal1 40986 54672 40986 54672 0 _031_
rlabel metal1 38502 55250 38502 55250 0 _032_
rlabel metal1 38364 56270 38364 56270 0 _033_
rlabel metal1 38318 55284 38318 55284 0 _034_
rlabel metal1 38042 55930 38042 55930 0 _035_
rlabel metal1 37398 55624 37398 55624 0 _036_
rlabel metal2 35558 56100 35558 56100 0 _037_
rlabel metal1 36570 56882 36570 56882 0 _038_
rlabel metal1 35282 56474 35282 56474 0 _039_
rlabel metal2 33626 56882 33626 56882 0 _040_
rlabel metal2 31786 56508 31786 56508 0 _041_
rlabel metal1 31372 56474 31372 56474 0 _042_
rlabel metal1 24058 57358 24058 57358 0 _043_
rlabel metal2 36478 56644 36478 56644 0 _044_
rlabel metal1 40434 56848 40434 56848 0 _045_
rlabel metal1 40388 57018 40388 57018 0 _046_
rlabel metal1 40020 57562 40020 57562 0 _047_
rlabel metal2 24058 55420 24058 55420 0 _048_
rlabel metal1 23598 56338 23598 56338 0 _049_
rlabel metal2 32430 53958 32430 53958 0 _050_
rlabel metal1 33028 54298 33028 54298 0 _051_
rlabel metal1 33948 56338 33948 56338 0 _052_
rlabel metal2 33074 55930 33074 55930 0 _053_
rlabel metal1 25438 55658 25438 55658 0 _054_
rlabel metal2 41630 54604 41630 54604 0 _055_
rlabel metal1 41492 54298 41492 54298 0 _056_
rlabel metal1 42458 55930 42458 55930 0 _057_
rlabel metal1 41630 56338 41630 56338 0 _058_
rlabel via2 41078 56355 41078 56355 0 _059_
rlabel metal2 25714 55692 25714 55692 0 _060_
rlabel metal1 24932 55726 24932 55726 0 _061_
rlabel metal1 31602 55658 31602 55658 0 _062_
rlabel metal2 31326 55556 31326 55556 0 _063_
rlabel metal1 30728 54570 30728 54570 0 _064_
rlabel metal2 30774 55522 30774 55522 0 _065_
rlabel metal2 30866 55284 30866 55284 0 _066_
rlabel metal1 26910 55794 26910 55794 0 _067_
rlabel metal1 40158 56270 40158 56270 0 _068_
rlabel metal1 40066 56372 40066 56372 0 _069_
rlabel metal2 39974 55522 39974 55522 0 _070_
rlabel metal2 40894 56134 40894 56134 0 _071_
rlabel metal1 40292 55386 40292 55386 0 _072_
rlabel metal2 39882 55981 39882 55981 0 _073_
rlabel metal2 26450 55964 26450 55964 0 _074_
rlabel metal1 26404 55726 26404 55726 0 _075_
rlabel metal2 28566 54468 28566 54468 0 _076_
rlabel metal2 28474 54570 28474 54570 0 _077_
rlabel metal1 29486 56882 29486 56882 0 _078_
rlabel metal1 29118 56372 29118 56372 0 _079_
rlabel metal1 29670 56780 29670 56780 0 _080_
rlabel metal2 29578 57188 29578 57188 0 _081_
rlabel metal1 28382 56202 28382 56202 0 _082_
rlabel metal1 37352 55386 37352 55386 0 _083_
rlabel metal2 36662 55964 36662 55964 0 _084_
rlabel metal2 36754 56134 36754 56134 0 _085_
rlabel metal1 43286 56882 43286 56882 0 _086_
rlabel metal1 36294 56780 36294 56780 0 _087_
rlabel metal1 29302 56236 29302 56236 0 _088_
rlabel metal1 24610 5746 24610 5746 0 _089_
rlabel metal2 36754 4352 36754 4352 0 _090_
rlabel metal1 26082 4114 26082 4114 0 _091_
rlabel metal1 25346 4182 25346 4182 0 _092_
rlabel metal2 25530 5406 25530 5406 0 _093_
rlabel metal1 25070 4522 25070 4522 0 _094_
rlabel metal1 24564 3570 24564 3570 0 _095_
rlabel metal1 23092 3434 23092 3434 0 _096_
rlabel metal1 24886 2346 24886 2346 0 _097_
rlabel metal1 26496 5746 26496 5746 0 _098_
rlabel metal1 27830 5338 27830 5338 0 _099_
rlabel metal2 27830 6494 27830 6494 0 _100_
rlabel metal2 25438 3774 25438 3774 0 _101_
rlabel metal2 24702 3536 24702 3536 0 _102_
rlabel metal1 26082 4012 26082 4012 0 _103_
rlabel metal1 24610 3094 24610 3094 0 _104_
rlabel metal1 28658 2312 28658 2312 0 _105_
rlabel metal2 26082 3638 26082 3638 0 _106_
rlabel metal1 28750 5134 28750 5134 0 _107_
rlabel metal2 29486 6290 29486 6290 0 _108_
rlabel metal1 30176 8330 30176 8330 0 _109_
rlabel metal1 29808 4522 29808 4522 0 _110_
rlabel via2 24702 2941 24702 2941 0 _111_
rlabel metal2 30866 4488 30866 4488 0 _112_
rlabel metal1 31096 7718 31096 7718 0 _113_
rlabel metal2 30682 3298 30682 3298 0 _114_
rlabel metal2 33258 3230 33258 3230 0 _115_
rlabel metal2 33074 6052 33074 6052 0 _116_
rlabel metal1 33028 7174 33028 7174 0 _117_
rlabel metal1 34546 4182 34546 4182 0 _118_
rlabel metal1 36478 3094 36478 3094 0 _119_
rlabel metal1 36156 2346 36156 2346 0 _120_
rlabel metal2 34454 6188 34454 6188 0 _121_
rlabel metal1 36294 4522 36294 4522 0 _122_
rlabel metal2 37490 3026 37490 3026 0 _123_
rlabel metal1 34408 52054 34408 52054 0 _124_
rlabel metal2 3726 58388 3726 58388 0 io_active
rlabel metal1 27554 55692 27554 55692 0 io_in[18]
rlabel metal1 29486 57460 29486 57460 0 io_in[19]
rlabel metal1 32246 57426 32246 57426 0 io_in[20]
rlabel metal2 35650 57494 35650 57494 0 io_in[21]
rlabel metal1 34822 57426 34822 57426 0 io_in[22]
rlabel metal1 36340 57426 36340 57426 0 io_in[23]
rlabel metal1 37674 57426 37674 57426 0 io_in[24]
rlabel metal2 38732 56814 38732 56814 0 io_in[25]
rlabel metal1 40112 54162 40112 54162 0 io_in[26]
rlabel metal2 45218 57290 45218 57290 0 io_in[27]
rlabel metal1 42872 57426 42872 57426 0 io_in[28]
rlabel metal1 45816 55930 45816 55930 0 io_in[29]
rlabel metal1 45724 57494 45724 57494 0 io_in[30]
rlabel metal1 47012 57426 47012 57426 0 io_in[31]
rlabel metal1 48438 57426 48438 57426 0 io_in[32]
rlabel metal1 49772 57426 49772 57426 0 io_in[33]
rlabel metal1 51290 57426 51290 57426 0 io_in[34]
rlabel metal1 52578 57494 52578 57494 0 io_in[35]
rlabel metal1 54142 57426 54142 57426 0 io_in[36]
rlabel metal1 55430 57426 55430 57426 0 io_in[37]
rlabel metal1 5198 57562 5198 57562 0 io_out[0]
rlabel metal1 19044 57562 19044 57562 0 io_out[10]
rlabel metal1 20378 57562 20378 57562 0 io_out[11]
rlabel metal2 22034 58395 22034 58395 0 io_out[12]
rlabel metal1 23138 57562 23138 57562 0 io_out[13]
rlabel metal1 25024 57562 25024 57562 0 io_out[14]
rlabel metal1 25944 57562 25944 57562 0 io_out[15]
rlabel metal1 27646 57562 27646 57562 0 io_out[16]
rlabel metal1 28658 57562 28658 57562 0 io_out[17]
rlabel metal1 10718 57562 10718 57562 0 io_out[4]
rlabel metal1 12098 57562 12098 57562 0 io_out[5]
rlabel metal1 13478 57562 13478 57562 0 io_out[6]
rlabel metal1 14858 57562 14858 57562 0 io_out[7]
rlabel metal1 16238 57562 16238 57562 0 io_out[8]
rlabel metal1 17618 57562 17618 57562 0 io_out[9]
rlabel metal2 26174 1775 26174 1775 0 la_data_out[32]
rlabel metal2 26450 2710 26450 2710 0 la_data_out[33]
rlabel metal2 26726 2098 26726 2098 0 la_data_out[34]
rlabel metal2 27002 2064 27002 2064 0 la_data_out[35]
rlabel metal2 27278 1554 27278 1554 0 la_data_out[36]
rlabel metal2 27554 3254 27554 3254 0 la_data_out[37]
rlabel metal2 27830 2098 27830 2098 0 la_data_out[38]
rlabel metal2 28106 3492 28106 3492 0 la_data_out[39]
rlabel metal2 28382 2200 28382 2200 0 la_data_out[40]
rlabel metal2 28658 1860 28658 1860 0 la_data_out[41]
rlabel metal2 28934 2370 28934 2370 0 la_data_out[42]
rlabel metal2 29210 1792 29210 1792 0 la_data_out[43]
rlabel metal2 29486 1622 29486 1622 0 la_data_out[44]
rlabel metal2 29762 2404 29762 2404 0 la_data_out[45]
rlabel metal2 30038 1792 30038 1792 0 la_data_out[46]
rlabel metal2 30314 3798 30314 3798 0 la_data_out[47]
rlabel metal2 30590 3254 30590 3254 0 la_data_out[48]
rlabel metal2 30866 1503 30866 1503 0 la_data_out[49]
rlabel metal2 31142 1622 31142 1622 0 la_data_out[50]
rlabel metal2 31418 1894 31418 1894 0 la_data_out[51]
rlabel metal2 31694 2387 31694 2387 0 la_data_out[52]
rlabel metal2 31970 2166 31970 2166 0 la_data_out[53]
rlabel metal2 32246 1860 32246 1860 0 la_data_out[54]
rlabel metal2 32522 1979 32522 1979 0 la_data_out[55]
rlabel metal2 32798 1792 32798 1792 0 la_data_out[56]
rlabel metal2 33074 2404 33074 2404 0 la_data_out[57]
rlabel metal2 33350 1826 33350 1826 0 la_data_out[58]
rlabel metal2 33626 1554 33626 1554 0 la_data_out[59]
rlabel metal2 33902 3288 33902 3288 0 la_data_out[60]
rlabel metal2 34178 2642 34178 2642 0 la_data_out[61]
rlabel metal2 34454 2166 34454 2166 0 la_data_out[62]
rlabel metal2 34730 3831 34730 3831 0 la_data_out[63]
rlabel metal2 5382 56712 5382 56712 0 net1
rlabel metal1 40572 55046 40572 55046 0 net10
rlabel metal2 35834 1826 35834 1826 0 net100
rlabel metal2 36110 2234 36110 2234 0 net101
rlabel metal2 36386 1520 36386 1520 0 net102
rlabel metal2 36662 1299 36662 1299 0 net103
rlabel metal2 36938 1792 36938 1792 0 net104
rlabel metal2 37214 2370 37214 2370 0 net105
rlabel metal2 37490 1299 37490 1299 0 net106
rlabel metal2 37766 1554 37766 1554 0 net107
rlabel metal2 38042 1894 38042 1894 0 net108
rlabel metal2 38318 1656 38318 1656 0 net109
rlabel metal1 42596 55726 42596 55726 0 net11
rlabel metal2 38594 2336 38594 2336 0 net110
rlabel metal2 38870 1826 38870 1826 0 net111
rlabel metal2 39146 1622 39146 1622 0 net112
rlabel metal2 39422 2132 39422 2132 0 net113
rlabel metal2 39698 1860 39698 1860 0 net114
rlabel metal2 39974 2200 39974 2200 0 net115
rlabel metal2 40250 1894 40250 1894 0 net116
rlabel metal2 40526 1554 40526 1554 0 net117
rlabel metal2 40802 2166 40802 2166 0 net118
rlabel metal2 41078 1826 41078 1826 0 net119
rlabel metal1 43194 56338 43194 56338 0 net12
rlabel metal2 41354 2132 41354 2132 0 net120
rlabel metal2 41630 1656 41630 1656 0 net121
rlabel metal2 41906 1792 41906 1792 0 net122
rlabel metal2 42182 1622 42182 1622 0 net123
rlabel metal2 42458 2132 42458 2132 0 net124
rlabel metal2 42734 1588 42734 1588 0 net125
rlabel metal2 43010 1826 43010 1826 0 net126
rlabel metal2 43286 2132 43286 2132 0 net127
rlabel metal2 43562 1792 43562 1792 0 net128
rlabel metal2 43838 1554 43838 1554 0 net129
rlabel metal2 40434 55760 40434 55760 0 net13
rlabel metal2 44114 2132 44114 2132 0 net130
rlabel metal2 44390 1826 44390 1826 0 net131
rlabel metal2 44666 1622 44666 1622 0 net132
rlabel metal2 44942 1792 44942 1792 0 net133
rlabel metal2 45218 1656 45218 1656 0 net134
rlabel metal2 45494 1860 45494 1860 0 net135
rlabel metal2 45770 1588 45770 1588 0 net136
rlabel metal2 46046 2132 46046 2132 0 net137
rlabel metal2 46322 1792 46322 1792 0 net138
rlabel metal2 46598 2132 46598 2132 0 net139
rlabel metal2 44942 56474 44942 56474 0 net14
rlabel metal2 46874 1860 46874 1860 0 net140
rlabel metal2 47150 1622 47150 1622 0 net141
rlabel metal2 47426 1554 47426 1554 0 net142
rlabel metal2 47702 1826 47702 1826 0 net143
rlabel metal2 47978 1690 47978 1690 0 net144
rlabel metal2 48254 2132 48254 2132 0 net145
rlabel metal2 48530 1792 48530 1792 0 net146
rlabel metal2 48806 1656 48806 1656 0 net147
rlabel metal2 49082 1826 49082 1826 0 net148
rlabel metal2 49358 2132 49358 2132 0 net149
rlabel metal2 45034 56610 45034 56610 0 net15
rlabel metal2 49634 1792 49634 1792 0 net150
rlabel metal2 49910 1622 49910 1622 0 net151
rlabel metal2 50186 2132 50186 2132 0 net152
rlabel metal2 50462 1095 50462 1095 0 net153
rlabel metal2 50738 1656 50738 1656 0 net154
rlabel metal2 51014 1826 51014 1826 0 net155
rlabel metal2 51290 1554 51290 1554 0 net156
rlabel metal2 51566 1792 51566 1792 0 net157
rlabel metal2 51842 1622 51842 1622 0 net158
rlabel metal2 52118 2132 52118 2132 0 net159
rlabel metal1 44850 55760 44850 55760 0 net16
rlabel metal2 52394 1826 52394 1826 0 net160
rlabel metal2 7682 1792 7682 1792 0 net161
rlabel metal2 8234 1588 8234 1588 0 net162
rlabel metal2 8602 1792 8602 1792 0 net163
rlabel metal2 8970 1588 8970 1588 0 net164
rlabel metal2 9338 2132 9338 2132 0 net165
rlabel metal2 9706 1656 9706 1656 0 net166
rlabel metal2 9982 1792 9982 1792 0 net167
rlabel metal2 10258 1588 10258 1588 0 net168
rlabel metal2 10534 1792 10534 1792 0 net169
rlabel metal1 44114 56814 44114 56814 0 net17
rlabel metal2 10810 2132 10810 2132 0 net170
rlabel metal2 11086 1792 11086 1792 0 net171
rlabel metal2 11362 1656 11362 1656 0 net172
rlabel metal2 11638 1792 11638 1792 0 net173
rlabel metal2 11914 1588 11914 1588 0 net174
rlabel metal2 12190 1792 12190 1792 0 net175
rlabel metal2 12466 2132 12466 2132 0 net176
rlabel metal2 12742 1622 12742 1622 0 net177
rlabel metal2 13018 1792 13018 1792 0 net178
rlabel metal2 13294 1588 13294 1588 0 net179
rlabel metal2 51658 56457 51658 56457 0 net18
rlabel metal2 13570 2132 13570 2132 0 net180
rlabel metal2 13846 1792 13846 1792 0 net181
rlabel metal2 14122 1588 14122 1588 0 net182
rlabel metal2 14398 1792 14398 1792 0 net183
rlabel metal2 14674 2132 14674 2132 0 net184
rlabel metal2 14950 1656 14950 1656 0 net185
rlabel metal2 15226 1792 15226 1792 0 net186
rlabel metal2 15502 2132 15502 2132 0 net187
rlabel metal2 15778 1554 15778 1554 0 net188
rlabel metal2 16054 1792 16054 1792 0 net189
rlabel metal2 52762 56253 52762 56253 0 net19
rlabel metal2 16330 1588 16330 1588 0 net190
rlabel metal2 16606 2132 16606 2132 0 net191
rlabel metal2 16882 1860 16882 1860 0 net192
rlabel metal2 17158 1792 17158 1792 0 net193
rlabel metal2 25346 5644 25346 5644 0 net194
rlabel metal2 25898 4828 25898 4828 0 net195
rlabel metal2 25898 3774 25898 3774 0 net196
rlabel metal1 23046 2618 23046 2618 0 net197
rlabel metal1 24334 2482 24334 2482 0 net198
rlabel metal1 25668 5678 25668 5678 0 net199
rlabel metal2 31878 55590 31878 55590 0 net2
rlabel metal1 45539 56338 45539 56338 0 net20
rlabel metal1 27002 6154 27002 6154 0 net200
rlabel metal2 27646 6528 27646 6528 0 net201
rlabel metal2 27278 4114 27278 4114 0 net202
rlabel metal2 27922 3910 27922 3910 0 net203
rlabel metal2 22862 3366 22862 3366 0 net204
rlabel metal1 24702 2618 24702 2618 0 net205
rlabel metal1 27370 2958 27370 2958 0 net206
rlabel metal1 28750 4114 28750 4114 0 net207
rlabel metal2 28934 5440 28934 5440 0 net208
rlabel metal1 29118 6834 29118 6834 0 net209
rlabel metal2 55430 56542 55430 56542 0 net21
rlabel metal1 30084 7854 30084 7854 0 net210
rlabel metal1 30084 4590 30084 4590 0 net211
rlabel metal2 36202 2652 36202 2652 0 net212
rlabel metal2 31326 4624 31326 4624 0 net213
rlabel metal1 31188 6698 31188 6698 0 net214
rlabel metal2 31510 3740 31510 3740 0 net215
rlabel metal2 33442 3468 33442 3468 0 net216
rlabel metal2 32522 6018 32522 6018 0 net217
rlabel metal1 33212 4794 33212 4794 0 net218
rlabel metal2 34546 4352 34546 4352 0 net219
rlabel metal2 5474 57052 5474 57052 0 net22
rlabel metal2 35742 3468 35742 3468 0 net220
rlabel metal2 36570 3026 36570 3026 0 net221
rlabel metal2 34270 5916 34270 5916 0 net222
rlabel metal2 36110 4828 36110 4828 0 net223
rlabel metal1 36708 3570 36708 3570 0 net224
rlabel metal1 34178 51578 34178 51578 0 net225
rlabel metal1 4692 57018 4692 57018 0 net226
rlabel metal1 5980 57426 5980 57426 0 net227
rlabel metal1 7360 57426 7360 57426 0 net228
rlabel metal1 8740 57426 8740 57426 0 net229
rlabel metal1 20838 57324 20838 57324 0 net23
rlabel metal1 10258 57018 10258 57018 0 net230
rlabel metal1 11500 57426 11500 57426 0 net231
rlabel metal1 12972 57018 12972 57018 0 net232
rlabel metal1 14260 57426 14260 57426 0 net233
rlabel metal1 16008 57018 16008 57018 0 net234
rlabel metal1 17020 57426 17020 57426 0 net235
rlabel metal1 18400 57426 18400 57426 0 net236
rlabel metal1 19964 57018 19964 57018 0 net237
rlabel metal1 21252 57018 21252 57018 0 net238
rlabel metal1 22632 56338 22632 56338 0 net239
rlabel metal2 20654 57324 20654 57324 0 net24
rlabel metal2 21482 57375 21482 57375 0 net240
rlabel metal1 24150 56950 24150 56950 0 net241
rlabel metal1 26772 54842 26772 54842 0 net242
rlabel metal1 27922 54842 27922 54842 0 net243
rlabel metal1 29854 54842 29854 54842 0 net244
rlabel metal1 30912 57426 30912 57426 0 net245
rlabel metal1 32338 56338 32338 56338 0 net246
rlabel metal1 34776 55930 34776 55930 0 net247
rlabel metal1 35604 54842 35604 54842 0 net248
rlabel metal1 36432 54842 36432 54842 0 net249
rlabel metal2 26266 56491 26266 56491 0 net25
rlabel metal1 37812 54842 37812 54842 0 net250
rlabel metal2 39146 57861 39146 57861 0 net251
rlabel metal2 40618 56627 40618 56627 0 net252
rlabel metal1 42228 55182 42228 55182 0 net253
rlabel metal2 46414 56848 46414 56848 0 net254
rlabel metal1 46138 56168 46138 56168 0 net255
rlabel metal1 46782 56950 46782 56950 0 net256
rlabel metal1 47794 57018 47794 57018 0 net257
rlabel metal1 49128 57018 49128 57018 0 net258
rlabel metal2 36110 56593 36110 56593 0 net26
rlabel metal1 23828 57018 23828 57018 0 net27
rlabel metal2 25622 56372 25622 56372 0 net28
rlabel metal2 26358 56780 26358 56780 0 net29
rlabel metal1 34362 56304 34362 56304 0 net3
rlabel metal2 29118 57222 29118 57222 0 net30
rlabel metal2 10994 57188 10994 57188 0 net31
rlabel metal2 12374 57630 12374 57630 0 net32
rlabel metal1 21390 57460 21390 57460 0 net33
rlabel metal2 15134 57664 15134 57664 0 net34
rlabel metal2 16514 57154 16514 57154 0 net35
rlabel metal2 17894 56916 17894 56916 0 net36
rlabel metal1 50462 57018 50462 57018 0 net37
rlabel metal1 51888 57018 51888 57018 0 net38
rlabel metal1 53222 57426 53222 57426 0 net39
rlabel metal2 32706 54740 32706 54740 0 net4
rlabel metal1 54372 57018 54372 57018 0 net40
rlabel metal1 55890 57426 55890 57426 0 net41
rlabel metal1 6532 57426 6532 57426 0 net42
rlabel metal1 7912 57426 7912 57426 0 net43
rlabel metal1 9292 57426 9292 57426 0 net44
rlabel metal1 29992 56338 29992 56338 0 net45
rlabel metal1 30820 57358 30820 57358 0 net46
rlabel metal1 33488 57018 33488 57018 0 net47
rlabel metal1 35006 54842 35006 54842 0 net48
rlabel metal1 37306 55250 37306 55250 0 net49
rlabel metal2 33028 56814 33028 56814 0 net5
rlabel metal2 41078 56848 41078 56848 0 net50
rlabel metal1 38272 54162 38272 54162 0 net51
rlabel metal2 39606 57725 39606 57725 0 net52
rlabel metal2 40986 57538 40986 57538 0 net53
rlabel metal1 43286 55216 43286 55216 0 net54
rlabel metal2 46230 56610 46230 56610 0 net55
rlabel metal1 45954 56270 45954 56270 0 net56
rlabel metal1 46966 56338 46966 56338 0 net57
rlabel metal1 48346 56882 48346 56882 0 net58
rlabel metal1 49680 56950 49680 56950 0 net59
rlabel metal1 35512 55114 35512 55114 0 net6
rlabel metal2 50646 58082 50646 58082 0 net60
rlabel metal1 52440 56950 52440 56950 0 net61
rlabel metal1 53452 57018 53452 57018 0 net62
rlabel metal1 54924 57018 54924 57018 0 net63
rlabel metal1 56212 57018 56212 57018 0 net64
rlabel metal2 17342 2132 17342 2132 0 net65
rlabel metal2 17618 1622 17618 1622 0 net66
rlabel metal2 17894 1792 17894 1792 0 net67
rlabel metal2 18170 2132 18170 2132 0 net68
rlabel metal2 18446 1656 18446 1656 0 net69
rlabel metal2 34638 56848 34638 56848 0 net7
rlabel metal2 18722 1792 18722 1792 0 net70
rlabel metal2 18998 2132 18998 2132 0 net71
rlabel metal2 19274 1622 19274 1622 0 net72
rlabel metal2 19550 1095 19550 1095 0 net73
rlabel metal2 19826 1367 19826 1367 0 net74
rlabel metal2 20102 1656 20102 1656 0 net75
rlabel metal2 20378 2132 20378 2132 0 net76
rlabel metal2 20654 2336 20654 2336 0 net77
rlabel metal2 20930 2132 20930 2132 0 net78
rlabel metal2 21206 1860 21206 1860 0 net79
rlabel metal2 35190 55318 35190 55318 0 net8
rlabel metal2 21482 2676 21482 2676 0 net80
rlabel metal2 21758 1826 21758 1826 0 net81
rlabel metal2 22034 2336 22034 2336 0 net82
rlabel metal2 22310 2200 22310 2200 0 net83
rlabel metal2 22586 2676 22586 2676 0 net84
rlabel metal2 22862 1622 22862 1622 0 net85
rlabel metal2 23138 2880 23138 2880 0 net86
rlabel metal2 23414 1860 23414 1860 0 net87
rlabel metal2 23690 2370 23690 2370 0 net88
rlabel metal2 23966 2744 23966 2744 0 net89
rlabel metal1 35604 55726 35604 55726 0 net9
rlabel metal2 24242 959 24242 959 0 net90
rlabel metal2 24518 1078 24518 1078 0 net91
rlabel metal2 24794 2948 24794 2948 0 net92
rlabel metal2 25070 1656 25070 1656 0 net93
rlabel metal2 25346 2200 25346 2200 0 net94
rlabel metal2 25622 1095 25622 1095 0 net95
rlabel metal2 25898 1418 25898 1418 0 net96
rlabel metal2 35006 1656 35006 1656 0 net97
rlabel metal2 35282 1163 35282 1163 0 net98
rlabel metal2 38686 2703 38686 2703 0 net99
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
