* NGSPICE file created from macro_decap_3.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_4 abstract view
.subckt sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_8 abstract view
.subckt sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

.subckt macro_decap_3 io_active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101]
+ la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108]
+ la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114]
+ la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120]
+ la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69]
+ la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81]
+ la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88]
+ la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94]
+ la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] vccd1 vssd1
+ wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__274__B1 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_294_ _044_ _085_ _087_ _124_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__a211oi_2
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_277_ _074_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XANTENNA__213__A_N net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_538__213 vssd1 vssd1 vccd1 vccd1 _538__213/HI net213 sky130_fd_sc_hd__conb_1
XFILLER_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_200_ net7 _000_ net6 vssd1 vssd1 vccd1 vccd1 _007_ sky130_fd_sc_hd__nand3b_1
XFILLER_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xmacro_decap_3_232 vssd1 vssd1 vccd1 vccd1 macro_decap_3_232/HI io_oeb[6] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_254 vssd1 vssd1 vccd1 vccd1 macro_decap_3_254/HI io_oeb[28] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_243 vssd1 vssd1 vccd1 vccd1 macro_decap_3_243/HI io_oeb[17] sky130_fd_sc_hd__conb_1
XFILLER_83_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input18_A io_in[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xmacro_decap_3_45 vssd1 vssd1 vccd1 vccd1 macro_decap_3_45/HI io_out[18] sky130_fd_sc_hd__conb_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_56 vssd1 vssd1 vccd1 vccd1 macro_decap_3_56/HI io_out[29] sky130_fd_sc_hd__conb_1
XFILLER_85_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmacro_decap_3_67 vssd1 vssd1 vccd1 vccd1 macro_decap_3_67/HI la_data_out[2] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_78 vssd1 vssd1 vccd1 vccd1 macro_decap_3_78/HI la_data_out[13] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_89 vssd1 vssd1 vccd1 vccd1 macro_decap_3_89/HI la_data_out[24] sky130_fd_sc_hd__conb_1
XFILLER_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_2
XFILLER_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_293_ _044_ _085_ _087_ vssd1 vssd1 vccd1 vccd1 _088_ sky130_fd_sc_hd__a21o_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_276_ net1 _073_ vssd1 vssd1 vccd1 vccd1 _074_ sky130_fd_sc_hd__and2_1
XFILLER_5_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_259_ _089_ _059_ vssd1 vssd1 vccd1 vccd1 _060_ sky130_fd_sc_hd__and2_1
XFILLER_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_233 vssd1 vssd1 vccd1 vccd1 macro_decap_3_233/HI io_oeb[7] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_244 vssd1 vssd1 vccd1 vccd1 macro_decap_3_244/HI io_oeb[18] sky130_fd_sc_hd__conb_1
XFILLER_16_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_255 vssd1 vssd1 vccd1 vccd1 macro_decap_3_255/HI io_oeb[29] sky130_fd_sc_hd__conb_1
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output31_A net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_523__198 vssd1 vssd1 vccd1 vccd1 _523__198/HI net198 sky130_fd_sc_hd__conb_1
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__295__C1 _089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmacro_decap_3_57 vssd1 vssd1 vccd1 vccd1 macro_decap_3_57/HI io_out[30] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_46 vssd1 vssd1 vccd1 vccd1 macro_decap_3_46/HI io_out[19] sky130_fd_sc_hd__conb_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmacro_decap_3_68 vssd1 vssd1 vccd1 vccd1 macro_decap_3_68/HI la_data_out[3] sky130_fd_sc_hd__conb_1
XFILLER_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_79 vssd1 vssd1 vccd1 vccd1 macro_decap_3_79/HI la_data_out[14] sky130_fd_sc_hd__conb_1
XFILLER_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_292_ net17 net20 _044_ _086_ vssd1 vssd1 vccd1 vccd1 _087_ sky130_fd_sc_hd__a211oi_2
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_275_ net21 _068_ _069_ _071_ _072_ vssd1 vssd1 vccd1 vccd1 _073_ sky130_fd_sc_hd__a32o_1
XFILLER_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_258_ net21 _056_ _058_ vssd1 vssd1 vccd1 vccd1 _059_ sky130_fd_sc_hd__o21a_1
X_189_ _092_ vssd1 vssd1 vccd1 vccd1 _096_ sky130_fd_sc_hd__inv_2
XFILLER_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xmacro_decap_3_245 vssd1 vssd1 vccd1 vccd1 macro_decap_3_245/HI io_oeb[19] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_234 vssd1 vssd1 vccd1 vccd1 macro_decap_3_234/HI io_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_16_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_256 vssd1 vssd1 vccd1 vccd1 macro_decap_3_256/HI io_oeb[30] sky130_fd_sc_hd__conb_1
XFILLER_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__236__A net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_528__203 vssd1 vssd1 vccd1 vccd1 _528__203/HI net203 sky130_fd_sc_hd__conb_1
XFILLER_81_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmacro_decap_3_58 vssd1 vssd1 vccd1 vccd1 macro_decap_3_58/HI io_out[31] sky130_fd_sc_hd__conb_1
XFILLER_97_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xmacro_decap_3_47 vssd1 vssd1 vccd1 vccd1 macro_decap_3_47/HI io_out[20] sky130_fd_sc_hd__conb_1
XFILLER_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmacro_decap_3_69 vssd1 vssd1 vccd1 vccd1 macro_decap_3_69/HI la_data_out[4] sky130_fd_sc_hd__conb_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_2
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_2
XFILLER_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__268__B1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_291_ net17 net20 net13 vssd1 vssd1 vccd1 vccd1 _086_ sky130_fd_sc_hd__o21a_1
XFILLER_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__244__A _089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_274_ _070_ _032_ net21 vssd1 vssd1 vccd1 vccd1 _072_ sky130_fd_sc_hd__a21oi_1
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_257_ net15 net20 _044_ _057_ vssd1 vssd1 vccd1 vccd1 _058_ sky130_fd_sc_hd__a211o_1
X_188_ _092_ vssd1 vssd1 vccd1 vccd1 _097_ sky130_fd_sc_hd__inv_2
XFILLER_6_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_235 vssd1 vssd1 vccd1 vccd1 macro_decap_3_235/HI io_oeb[9] sky130_fd_sc_hd__conb_1
XFILLER_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_257 vssd1 vssd1 vccd1 vccd1 macro_decap_3_257/HI io_oeb[31] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_246 vssd1 vssd1 vccd1 vccd1 macro_decap_3_246/HI io_oeb[20] sky130_fd_sc_hd__conb_1
XFILLER_34_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__295__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__157__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmacro_decap_3_37 vssd1 vssd1 vccd1 vccd1 macro_decap_3_37/HI io_oeb[33] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_59 vssd1 vssd1 vccd1 vccd1 macro_decap_3_59/HI io_out[32] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_48 vssd1 vssd1 vccd1 vccd1 macro_decap_3_48/HI io_out[21] sky130_fd_sc_hd__conb_1
XFILLER_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_2
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input16_A io_in[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input8_A io_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_290_ _083_ _084_ vssd1 vssd1 vccd1 vccd1 _085_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__170__A _089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_273_ _070_ _032_ vssd1 vssd1 vccd1 vccd1 _071_ sky130_fd_sc_hd__or2_1
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_519__194 vssd1 vssd1 vccd1 vccd1 _519__194/HI net194 sky130_fd_sc_hd__conb_1
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_256_ net15 net20 net11 vssd1 vssd1 vccd1 vccd1 _057_ sky130_fd_sc_hd__o21a_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_187_ _092_ vssd1 vssd1 vccd1 vccd1 _098_ sky130_fd_sc_hd__inv_2
XFILLER_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_236 vssd1 vssd1 vccd1 vccd1 macro_decap_3_236/HI io_oeb[10] sky130_fd_sc_hd__conb_1
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmacro_decap_3_258 vssd1 vssd1 vccd1 vccd1 macro_decap_3_258/HI io_oeb[32] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_247 vssd1 vssd1 vccd1 vccd1 macro_decap_3_247/HI io_oeb[21] sky130_fd_sc_hd__conb_1
XFILLER_70_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_239_ net6 net19 net2 _042_ vssd1 vssd1 vccd1 vccd1 _043_ sky130_fd_sc_hd__a31o_1
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__286__A2 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmacro_decap_3_38 vssd1 vssd1 vccd1 vccd1 macro_decap_3_38/HI io_oeb[34] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_49 vssd1 vssd1 vccd1 vccd1 macro_decap_3_49/HI io_out[22] sky130_fd_sc_hd__conb_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_2
Xoutput35 net35 vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__buf_2
XFILLER_88_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_272_ net12 _025_ vssd1 vssd1 vccd1 vccd1 _070_ sky130_fd_sc_hd__xor2_1
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_539_ net214 _113_ vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__ebufn_8
XFILLER_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__181__A _089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_255_ _055_ _030_ vssd1 vssd1 vccd1 vccd1 _056_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_186_ _092_ vssd1 vssd1 vccd1 vccd1 _099_ sky130_fd_sc_hd__inv_2
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_226 vssd1 vssd1 vccd1 vccd1 macro_decap_3_226/HI io_oeb[0] sky130_fd_sc_hd__conb_1
XFILLER_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_248 vssd1 vssd1 vccd1 vccd1 macro_decap_3_248/HI io_oeb[22] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_237 vssd1 vssd1 vccd1 vccd1 macro_decap_3_237/HI io_oeb[11] sky130_fd_sc_hd__conb_1
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__231__B1 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_238_ net6 net2 _041_ vssd1 vssd1 vccd1 vccd1 _042_ sky130_fd_sc_hd__o21a_1
X_169_ _090_ vssd1 vssd1 vccd1 vccd1 _114_ sky130_fd_sc_hd__inv_2
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_output22_A net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmacro_decap_3_39 vssd1 vssd1 vccd1 vccd1 macro_decap_3_39/HI io_oeb[35] sky130_fd_sc_hd__conb_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_2
Xoutput36 net36 vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__buf_2
XFILLER_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input21_A io_in[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_271_ net20 net12 vssd1 vssd1 vccd1 vccd1 _069_ sky130_fd_sc_hd__or2_1
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_538_ net213 _112_ vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__ebufn_8
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_254_ _031_ _029_ vssd1 vssd1 vccd1 vccd1 _055_ sky130_fd_sc_hd__or2b_1
XFILLER_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_185_ _092_ vssd1 vssd1 vccd1 vccd1 _100_ sky130_fd_sc_hd__inv_2
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__192__A _089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_227 vssd1 vssd1 vccd1 vccd1 macro_decap_3_227/HI io_oeb[1] sky130_fd_sc_hd__conb_1
XFILLER_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_238 vssd1 vssd1 vccd1 vccd1 macro_decap_3_238/HI io_oeb[12] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_249 vssd1 vssd1 vccd1 vccd1 macro_decap_3_249/HI io_oeb[23] sky130_fd_sc_hd__conb_1
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_237_ net6 net2 _040_ net18 vssd1 vssd1 vccd1 vccd1 _041_ sky130_fd_sc_hd__o2bb2a_1
X_168_ _090_ vssd1 vssd1 vccd1 vccd1 _115_ sky130_fd_sc_hd__inv_2
XFILLER_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input14_A io_in[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input6_A io_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_270_ net20 net12 net16 vssd1 vssd1 vccd1 vccd1 _068_ sky130_fd_sc_hd__a21o_1
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_537_ net212 _111_ vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__ebufn_8
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_253_ net19 _051_ _053_ vssd1 vssd1 vccd1 vccd1 _054_ sky130_fd_sc_hd__o21a_1
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_184_ _092_ vssd1 vssd1 vccd1 vccd1 _101_ sky130_fd_sc_hd__inv_2
XFILLER_89_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_228 vssd1 vssd1 vccd1 vccd1 macro_decap_3_228/HI io_oeb[2] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_239 vssd1 vssd1 vccd1 vccd1 macro_decap_3_239/HI io_oeb[13] sky130_fd_sc_hd__conb_1
XFILLER_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_236_ net19 vssd1 vssd1 vccd1 vccd1 _040_ sky130_fd_sc_hd__inv_2
XFILLER_10_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_167_ _090_ vssd1 vssd1 vccd1 vccd1 _116_ sky130_fd_sc_hd__inv_2
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_541__216 vssd1 vssd1 vccd1 vccd1 _541__216/HI net216 sky130_fd_sc_hd__conb_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_219_ net12 _025_ vssd1 vssd1 vccd1 vccd1 _026_ sky130_fd_sc_hd__or2_1
XFILLER_97_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_2
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_547__222 vssd1 vssd1 vccd1 vccd1 _547__222/HI net222 sky130_fd_sc_hd__conb_1
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_536_ net211 _110_ vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__ebufn_8
XFILLER_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_252_ net7 net18 _040_ _052_ vssd1 vssd1 vccd1 vccd1 _053_ sky130_fd_sc_hd__a211o_1
XFILLER_80_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_183_ _092_ vssd1 vssd1 vccd1 vccd1 _102_ sky130_fd_sc_hd__inv_2
XFILLER_89_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_519_ net194 _093_ vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__ebufn_8
XFILLER_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmacro_decap_3_229 vssd1 vssd1 vccd1 vccd1 macro_decap_3_229/HI io_oeb[3] sky130_fd_sc_hd__conb_1
XFILLER_83_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_235_ _019_ _039_ net31 net32 vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__o22a_1
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_166_ _090_ vssd1 vssd1 vccd1 vccd1 _117_ sky130_fd_sc_hd__inv_2
XFILLER_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_218_ net16 _024_ vssd1 vssd1 vccd1 vccd1 _025_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_2
XFILLER_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_535_ net210 _109_ vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__ebufn_8
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_251_ net7 net18 net3 vssd1 vssd1 vccd1 vccd1 _052_ sky130_fd_sc_hd__o21a_1
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_182_ _092_ vssd1 vssd1 vccd1 vccd1 _103_ sky130_fd_sc_hd__inv_2
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_234_ _124_ _017_ _018_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__nor3_1
XFILLER_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_165_ _090_ vssd1 vssd1 vccd1 vccd1 _118_ sky130_fd_sc_hd__inv_2
XFILLER_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_217_ net14 net15 _020_ vssd1 vssd1 vccd1 vccd1 _024_ sky130_fd_sc_hd__o21a_1
XFILLER_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_2
XFILLER_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_531__206 vssd1 vssd1 vccd1 vccd1 _531__206/HI net206 sky130_fd_sc_hd__conb_1
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input12_A io_in[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_534_ net209 _108_ vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__ebufn_8
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__252__A2 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input4_A io_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__243__A2 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_250_ _050_ _010_ vssd1 vssd1 vccd1 vccd1 _051_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_181_ _089_ vssd1 vssd1 vccd1 vccd1 _092_ sky130_fd_sc_hd__buf_4
XFILLER_22_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_537__212 vssd1 vssd1 vccd1 vccd1 _537__212/HI net212 sky130_fd_sc_hd__conb_1
XFILLER_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_233_ _124_ _037_ _038_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__nor3_2
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_164_ _090_ vssd1 vssd1 vccd1 vccd1 _119_ sky130_fd_sc_hd__inv_2
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_216_ net13 _022_ vssd1 vssd1 vccd1 vccd1 _023_ sky130_fd_sc_hd__or2_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_550_ net225 _124_ vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__ebufn_8
XFILLER_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_533_ net208 _107_ vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__ebufn_8
XFILLER_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_180_ _091_ vssd1 vssd1 vccd1 vccd1 _104_ sky130_fd_sc_hd__inv_2
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_232_ _037_ _038_ vssd1 vssd1 vccd1 vccd1 _039_ sky130_fd_sc_hd__or2_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_163_ _090_ vssd1 vssd1 vccd1 vccd1 _120_ sky130_fd_sc_hd__inv_2
XFILLER_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_215_ net17 _021_ vssd1 vssd1 vccd1 vccd1 _022_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_522__197 vssd1 vssd1 vccd1 vccd1 _522__197/HI net197 sky130_fd_sc_hd__conb_1
XFILLER_0_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__264__A1 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_190 vssd1 vssd1 vccd1 vccd1 macro_decap_3_190/HI wbs_dat_o[28] sky130_fd_sc_hd__conb_1
XFILLER_16_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_532_ net207 _106_ vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__ebufn_8
XFILLER_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__237__B2 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_231_ _036_ _023_ _035_ net21 vssd1 vssd1 vccd1 vccd1 _038_ sky130_fd_sc_hd__a31o_1
XFILLER_23_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_162_ _090_ vssd1 vssd1 vccd1 vccd1 _121_ sky130_fd_sc_hd__inv_2
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput1 io_active vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
XFILLER_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_527__202 vssd1 vssd1 vccd1 vccd1 _527__202/HI net202 sky130_fd_sc_hd__conb_1
XFILLER_45_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_214_ net16 net14 net15 _020_ vssd1 vssd1 vccd1 vccd1 _021_ sky130_fd_sc_hd__o31a_1
XFILLER_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_180 vssd1 vssd1 vccd1 vccd1 macro_decap_3_180/HI wbs_dat_o[18] sky130_fd_sc_hd__conb_1
XFILLER_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_191 vssd1 vssd1 vccd1 vccd1 macro_decap_3_191/HI wbs_dat_o[29] sky130_fd_sc_hd__conb_1
XFILLER_31_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_531_ net206 _105_ vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__ebufn_8
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input10_A io_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_544__219 vssd1 vssd1 vccd1 vccd1 _544__219/HI net219 sky130_fd_sc_hd__conb_1
XFILLER_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input2_A io_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_230_ _023_ _035_ _036_ vssd1 vssd1 vccd1 vccd1 _037_ sky130_fd_sc_hd__a21oi_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_161_ _090_ vssd1 vssd1 vccd1 vccd1 _122_ sky130_fd_sc_hd__inv_2
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput2 io_in[18] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_96_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_213_ net21 net20 vssd1 vssd1 vccd1 vccd1 _020_ sky130_fd_sc_hd__nand2b_1
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_181 vssd1 vssd1 vccd1 vccd1 macro_decap_3_181/HI wbs_dat_o[19] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_170 vssd1 vssd1 vccd1 vccd1 macro_decap_3_170/HI wbs_dat_o[8] sky130_fd_sc_hd__conb_1
XFILLER_16_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_192 vssd1 vssd1 vccd1 vccd1 macro_decap_3_192/HI wbs_dat_o[30] sky130_fd_sc_hd__conb_1
XFILLER_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_530_ net205 _104_ vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__ebufn_8
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_160_ _090_ vssd1 vssd1 vccd1 vccd1 _123_ sky130_fd_sc_hd__inv_2
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_289_ _033_ _023_ vssd1 vssd1 vccd1 vccd1 _084_ sky130_fd_sc_hd__and2b_1
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput3 io_in[19] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ _017_ _018_ vssd1 vssd1 vccd1 vccd1 _019_ sky130_fd_sc_hd__or2_1
XFILLER_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__258__A1 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xmacro_decap_3_171 vssd1 vssd1 vccd1 vccd1 macro_decap_3_171/HI wbs_dat_o[9] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_160 vssd1 vssd1 vccd1 vccd1 macro_decap_3_160/HI la_data_out[127] sky130_fd_sc_hd__conb_1
XFILLER_71_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_193 vssd1 vssd1 vccd1 vccd1 macro_decap_3_193/HI wbs_dat_o[31] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_182 vssd1 vssd1 vccd1 vccd1 macro_decap_3_182/HI wbs_dat_o[20] sky130_fd_sc_hd__conb_1
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_550__225 vssd1 vssd1 vccd1 vccd1 _550__225/HI net225 sky130_fd_sc_hd__conb_1
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_288_ _026_ _032_ _034_ vssd1 vssd1 vccd1 vccd1 _083_ sky130_fd_sc_hd__a21o_1
XFILLER_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput4 io_in[20] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_534__209 vssd1 vssd1 vccd1 vccd1 _534__209/HI net209 sky130_fd_sc_hd__conb_1
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_211_ _016_ _003_ _015_ net19 vssd1 vssd1 vccd1 vccd1 _018_ sky130_fd_sc_hd__a31o_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__285__A2 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__158__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_172 vssd1 vssd1 vccd1 vccd1 macro_decap_3_172/HI wbs_dat_o[10] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_161 vssd1 vssd1 vccd1 vccd1 macro_decap_3_161/HI wbs_ack_o sky130_fd_sc_hd__conb_1
Xmacro_decap_3_150 vssd1 vssd1 vccd1 vccd1 macro_decap_3_150/HI la_data_out[117] sky130_fd_sc_hd__conb_1
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_183 vssd1 vssd1 vccd1 vccd1 macro_decap_3_183/HI wbs_dat_o[21] sky130_fd_sc_hd__conb_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__261__A _089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_287_ _080_ _081_ vssd1 vssd1 vccd1 vccd1 _082_ sky130_fd_sc_hd__nor2_1
XFILLER_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput5 io_in[21] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_210_ _003_ _015_ _016_ vssd1 vssd1 vccd1 vccd1 _017_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input19_A io_in[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__259__A _089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xmacro_decap_3_162 vssd1 vssd1 vccd1 vccd1 macro_decap_3_162/HI wbs_dat_o[0] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_140 vssd1 vssd1 vccd1 vccd1 macro_decap_3_140/HI la_data_out[107] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_151 vssd1 vssd1 vccd1 vccd1 macro_decap_3_151/HI la_data_out[118] sky130_fd_sc_hd__conb_1
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_184 vssd1 vssd1 vccd1 vccd1 macro_decap_3_184/HI wbs_dat_o[22] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_173 vssd1 vssd1 vccd1 vccd1 macro_decap_3_173/HI wbs_dat_o[11] sky130_fd_sc_hd__conb_1
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_286_ net9 net18 _040_ vssd1 vssd1 vccd1 vccd1 _081_ sky130_fd_sc_hd__a21o_1
XFILLER_81_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput6 io_in[22] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_269_ net19 _062_ _063_ _065_ _066_ vssd1 vssd1 vccd1 vccd1 _067_ sky130_fd_sc_hd__a32o_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_540__215 vssd1 vssd1 vccd1 vccd1 _540__215/HI net215 sky130_fd_sc_hd__conb_1
XFILLER_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput20 io_in[36] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_2
XFILLER_69_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_141 vssd1 vssd1 vccd1 vccd1 macro_decap_3_141/HI la_data_out[108] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_163 vssd1 vssd1 vccd1 vccd1 macro_decap_3_163/HI wbs_dat_o[1] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_130 vssd1 vssd1 vccd1 vccd1 macro_decap_3_130/HI la_data_out[97] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_152 vssd1 vssd1 vccd1 vccd1 macro_decap_3_152/HI la_data_out[119] sky130_fd_sc_hd__conb_1
XFILLER_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_174 vssd1 vssd1 vccd1 vccd1 macro_decap_3_174/HI wbs_dat_o[12] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_185 vssd1 vssd1 vccd1 vccd1 macro_decap_3_185/HI wbs_dat_o[23] sky130_fd_sc_hd__conb_1
XFILLER_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_546__221 vssd1 vssd1 vccd1 vccd1 _546__221/HI net221 sky130_fd_sc_hd__conb_1
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_285_ net9 net18 net5 vssd1 vssd1 vccd1 vccd1 _080_ sky130_fd_sc_hd__o21a_1
XFILLER_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput7 io_in[23] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__278__A _089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_268_ _064_ _012_ net19 vssd1 vssd1 vccd1 vccd1 _066_ sky130_fd_sc_hd__a21oi_1
X_199_ net4 _005_ vssd1 vssd1 vccd1 vccd1 _006_ sky130_fd_sc_hd__or2_1
XFILLER_6_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput21 io_in[37] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_2
Xinput10 io_in[26] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_120 vssd1 vssd1 vccd1 vccd1 macro_decap_3_120/HI la_data_out[87] sky130_fd_sc_hd__conb_1
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmacro_decap_3_153 vssd1 vssd1 vccd1 vccd1 macro_decap_3_153/HI la_data_out[120] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_131 vssd1 vssd1 vccd1 vccd1 macro_decap_3_131/HI la_data_out[98] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_142 vssd1 vssd1 vccd1 vccd1 macro_decap_3_142/HI la_data_out[109] sky130_fd_sc_hd__conb_1
XFILLER_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xmacro_decap_3_186 vssd1 vssd1 vccd1 vccd1 macro_decap_3_186/HI wbs_dat_o[24] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_175 vssd1 vssd1 vccd1 vccd1 macro_decap_3_175/HI wbs_dat_o[13] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_164 vssd1 vssd1 vccd1 vccd1 macro_decap_3_164/HI wbs_dat_o[2] sky130_fd_sc_hd__conb_1
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__193__A_N net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_284_ net19 _078_ vssd1 vssd1 vccd1 vccd1 _079_ sky130_fd_sc_hd__nor2_1
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput8 io_in[24] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__193__B net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_267_ _064_ _012_ vssd1 vssd1 vccd1 vccd1 _065_ sky130_fd_sc_hd__or2_1
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_198_ net8 _004_ vssd1 vssd1 vccd1 vccd1 _005_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput11 io_in[27] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_110 vssd1 vssd1 vccd1 vccd1 macro_decap_3_110/HI la_data_out[77] sky130_fd_sc_hd__conb_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_121 vssd1 vssd1 vccd1 vccd1 macro_decap_3_121/HI la_data_out[88] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_132 vssd1 vssd1 vccd1 vccd1 macro_decap_3_132/HI la_data_out[99] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_143 vssd1 vssd1 vccd1 vccd1 macro_decap_3_143/HI la_data_out[110] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_154 vssd1 vssd1 vccd1 vccd1 macro_decap_3_154/HI la_data_out[121] sky130_fd_sc_hd__conb_1
XFILLER_16_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_187 vssd1 vssd1 vccd1 vccd1 macro_decap_3_187/HI wbs_dat_o[25] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_165 vssd1 vssd1 vccd1 vccd1 macro_decap_3_165/HI wbs_dat_o[3] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_176 vssd1 vssd1 vccd1 vccd1 macro_decap_3_176/HI wbs_dat_o[14] sky130_fd_sc_hd__conb_1
XFILLER_12_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_530__205 vssd1 vssd1 vccd1 vccd1 _530__205/HI net205 sky130_fd_sc_hd__conb_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input17_A io_in[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input9_A io_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_536__211 vssd1 vssd1 vccd1 vccd1 _536__211/HI net211 sky130_fd_sc_hd__conb_1
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_283_ _076_ _077_ vssd1 vssd1 vccd1 vccd1 _078_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput9 io_in[25] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_266_ net4 _005_ vssd1 vssd1 vccd1 vccd1 _064_ sky130_fd_sc_hd__xor2_1
X_197_ net6 net7 _000_ vssd1 vssd1 vccd1 vccd1 _004_ sky130_fd_sc_hd__o21a_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput12 io_in[28] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__dlymetal6s2s_1
X_249_ _011_ _009_ vssd1 vssd1 vccd1 vccd1 _050_ sky130_fd_sc_hd__or2b_1
XFILLER_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_100 vssd1 vssd1 vccd1 vccd1 macro_decap_3_100/HI la_data_out[67] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_111 vssd1 vssd1 vccd1 vccd1 macro_decap_3_111/HI la_data_out[78] sky130_fd_sc_hd__conb_1
XFILLER_16_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_144 vssd1 vssd1 vccd1 vccd1 macro_decap_3_144/HI la_data_out[111] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_122 vssd1 vssd1 vccd1 vccd1 macro_decap_3_122/HI la_data_out[89] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_133 vssd1 vssd1 vccd1 vccd1 macro_decap_3_133/HI la_data_out[100] sky130_fd_sc_hd__conb_1
XFILLER_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_155 vssd1 vssd1 vccd1 vccd1 macro_decap_3_155/HI la_data_out[122] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_177 vssd1 vssd1 vccd1 vccd1 macro_decap_3_177/HI wbs_dat_o[15] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_166 vssd1 vssd1 vccd1 vccd1 macro_decap_3_166/HI wbs_dat_o[4] sky130_fd_sc_hd__conb_1
XFILLER_43_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_188 vssd1 vssd1 vccd1 vccd1 macro_decap_3_188/HI wbs_dat_o[26] sky130_fd_sc_hd__conb_1
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__251__A2 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_282_ _013_ _003_ vssd1 vssd1 vccd1 vccd1 _077_ sky130_fd_sc_hd__and2b_1
XFILLER_41_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_549_ net224 _123_ vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__ebufn_8
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_265_ net18 net4 vssd1 vssd1 vccd1 vccd1 _063_ sky130_fd_sc_hd__or2_1
XFILLER_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_196_ net5 _002_ vssd1 vssd1 vccd1 vccd1 _003_ sky130_fd_sc_hd__or2_1
XFILLER_6_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_521__196 vssd1 vssd1 vccd1 vccd1 _521__196/HI net196 sky130_fd_sc_hd__conb_1
XFILLER_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput13 io_in[29] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_248_ _043_ _047_ net23 net27 vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_179_ _091_ vssd1 vssd1 vccd1 vccd1 _105_ sky130_fd_sc_hd__inv_2
XFILLER_6_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmacro_decap_3_101 vssd1 vssd1 vccd1 vccd1 macro_decap_3_101/HI la_data_out[68] sky130_fd_sc_hd__conb_1
XFILLER_83_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_134 vssd1 vssd1 vccd1 vccd1 macro_decap_3_134/HI la_data_out[101] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_112 vssd1 vssd1 vccd1 vccd1 macro_decap_3_112/HI la_data_out[79] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_123 vssd1 vssd1 vccd1 vccd1 macro_decap_3_123/HI la_data_out[90] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_145 vssd1 vssd1 vccd1 vccd1 macro_decap_3_145/HI la_data_out[112] sky130_fd_sc_hd__conb_1
XFILLER_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_178 vssd1 vssd1 vccd1 vccd1 macro_decap_3_178/HI wbs_dat_o[16] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_156 vssd1 vssd1 vccd1 vccd1 macro_decap_3_156/HI la_data_out[123] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_167 vssd1 vssd1 vccd1 vccd1 macro_decap_3_167/HI wbs_dat_o[5] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_189 vssd1 vssd1 vccd1 vccd1 macro_decap_3_189/HI wbs_dat_o[27] sky130_fd_sc_hd__conb_1
XFILLER_24_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_281_ _006_ _012_ _014_ vssd1 vssd1 vccd1 vccd1 _076_ sky130_fd_sc_hd__a21oi_1
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_548_ net223 _122_ vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__ebufn_8
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_526__201 vssd1 vssd1 vccd1 vccd1 _526__201/HI net201 sky130_fd_sc_hd__conb_1
XFILLER_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_264_ net18 net4 net8 vssd1 vssd1 vccd1 vccd1 _062_ sky130_fd_sc_hd__a21o_1
X_195_ net9 _001_ vssd1 vssd1 vccd1 vccd1 _002_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput14 io_in[30] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_2
X_247_ _049_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_178_ _091_ vssd1 vssd1 vccd1 vccd1 _106_ sky130_fd_sc_hd__inv_2
XFILLER_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_102 vssd1 vssd1 vccd1 vccd1 macro_decap_3_102/HI la_data_out[69] sky130_fd_sc_hd__conb_1
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_113 vssd1 vssd1 vccd1 vccd1 macro_decap_3_113/HI la_data_out[80] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_124 vssd1 vssd1 vccd1 vccd1 macro_decap_3_124/HI la_data_out[91] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_135 vssd1 vssd1 vccd1 vccd1 macro_decap_3_135/HI la_data_out[102] sky130_fd_sc_hd__conb_1
XFILLER_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmacro_decap_3_157 vssd1 vssd1 vccd1 vccd1 macro_decap_3_157/HI la_data_out[124] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_168 vssd1 vssd1 vccd1 vccd1 macro_decap_3_168/HI wbs_dat_o[6] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_146 vssd1 vssd1 vccd1 vccd1 macro_decap_3_146/HI la_data_out[113] sky130_fd_sc_hd__conb_1
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_179 vssd1 vssd1 vccd1 vccd1 macro_decap_3_179/HI wbs_dat_o[17] sky130_fd_sc_hd__conb_1
XFILLER_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input15_A io_in[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_543__218 vssd1 vssd1 vccd1 vccd1 _543__218/HI net218 sky130_fd_sc_hd__conb_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input7_A io_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_280_ _067_ _073_ net25 net29 vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__o2bb2a_1
XFILLER_14_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_547_ net222 _121_ vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__ebufn_8
XFILLER_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_263_ _054_ _059_ net24 net28 vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__o2bb2a_1
XFILLER_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_194_ net8 net6 net7 _000_ vssd1 vssd1 vccd1 vccd1 _001_ sky130_fd_sc_hd__o31a_1
XFILLER_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_549__224 vssd1 vssd1 vccd1 vccd1 _549__224/HI net224 sky130_fd_sc_hd__conb_1
XFILLER_28_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput15 io_in[31] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__dlymetal6s2s_1
X_246_ _089_ _043_ vssd1 vssd1 vccd1 vccd1 _049_ sky130_fd_sc_hd__and2_1
X_177_ _091_ vssd1 vssd1 vccd1 vccd1 _107_ sky130_fd_sc_hd__inv_2
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_136 vssd1 vssd1 vccd1 vccd1 macro_decap_3_136/HI la_data_out[103] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_103 vssd1 vssd1 vccd1 vccd1 macro_decap_3_103/HI la_data_out[70] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_114 vssd1 vssd1 vccd1 vccd1 macro_decap_3_114/HI la_data_out[81] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_125 vssd1 vssd1 vccd1 vccd1 macro_decap_3_125/HI la_data_out[92] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_169 vssd1 vssd1 vccd1 vccd1 macro_decap_3_169/HI wbs_dat_o[7] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_147 vssd1 vssd1 vccd1 vccd1 macro_decap_3_147/HI la_data_out[114] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_158 vssd1 vssd1 vccd1 vccd1 macro_decap_3_158/HI la_data_out[125] sky130_fd_sc_hd__conb_1
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_229_ net17 _020_ _021_ vssd1 vssd1 vccd1 vccd1 _036_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_546_ net221 _120_ vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__ebufn_8
XFILLER_17_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_262_ _061_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_193_ net19 net18 vssd1 vssd1 vccd1 vccd1 _000_ sky130_fd_sc_hd__nand2b_1
XFILLER_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_529_ net204 _103_ vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__ebufn_8
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_245_ _048_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput16 io_in[32] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_176_ _091_ vssd1 vssd1 vccd1 vccd1 _108_ sky130_fd_sc_hd__inv_2
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_126 vssd1 vssd1 vccd1 vccd1 macro_decap_3_126/HI la_data_out[93] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_115 vssd1 vssd1 vccd1 vccd1 macro_decap_3_115/HI la_data_out[82] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_104 vssd1 vssd1 vccd1 vccd1 macro_decap_3_104/HI la_data_out[71] sky130_fd_sc_hd__conb_1
XFILLER_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_148 vssd1 vssd1 vccd1 vccd1 macro_decap_3_148/HI la_data_out[115] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_137 vssd1 vssd1 vccd1 vccd1 macro_decap_3_137/HI la_data_out[104] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_159 vssd1 vssd1 vccd1 vccd1 macro_decap_3_159/HI la_data_out[126] sky130_fd_sc_hd__conb_1
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_228_ _026_ _032_ _033_ _034_ vssd1 vssd1 vccd1 vccd1 _035_ sky130_fd_sc_hd__a211o_1
X_159_ _089_ vssd1 vssd1 vccd1 vccd1 _090_ sky130_fd_sc_hd__buf_4
XFILLER_6_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input20_A io_in[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_545_ net220 _119_ vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__ebufn_8
XFILLER_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_261_ _089_ _054_ vssd1 vssd1 vccd1 vccd1 _061_ sky130_fd_sc_hd__and2_1
X_192_ _089_ vssd1 vssd1 vccd1 vccd1 _093_ sky130_fd_sc_hd__inv_2
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_533__208 vssd1 vssd1 vccd1 vccd1 _533__208/HI net208 sky130_fd_sc_hd__conb_1
XFILLER_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_528_ net203 _102_ vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__ebufn_8
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__275__A1 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_244_ _089_ _047_ vssd1 vssd1 vccd1 vccd1 _048_ sky130_fd_sc_hd__and2_1
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput17 io_in[33] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_175_ _091_ vssd1 vssd1 vccd1 vccd1 _109_ sky130_fd_sc_hd__inv_2
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_105 vssd1 vssd1 vccd1 vccd1 macro_decap_3_105/HI la_data_out[72] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_116 vssd1 vssd1 vccd1 vccd1 macro_decap_3_116/HI la_data_out[83] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_127 vssd1 vssd1 vccd1 vccd1 macro_decap_3_127/HI la_data_out[94] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_138 vssd1 vssd1 vccd1 vccd1 macro_decap_3_138/HI la_data_out[105] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_149 vssd1 vssd1 vccd1 vccd1 macro_decap_3_149/HI la_data_out[116] sky130_fd_sc_hd__conb_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__240__A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_539__214 vssd1 vssd1 vccd1 vccd1 _539__214/HI net214 sky130_fd_sc_hd__conb_1
X_227_ net12 _025_ vssd1 vssd1 vccd1 vccd1 _034_ sky130_fd_sc_hd__and2_1
X_158_ net1 vssd1 vssd1 vccd1 vccd1 _089_ sky130_fd_sc_hd__buf_4
XFILLER_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input13_A io_in[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_544_ net219 _118_ vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__ebufn_8
XFILLER_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input5_A io_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_260_ _060_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_191_ _092_ vssd1 vssd1 vccd1 vccd1 _094_ sky130_fd_sc_hd__inv_2
XFILLER_41_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_90 vssd1 vssd1 vccd1 vccd1 macro_decap_3_90/HI la_data_out[25] sky130_fd_sc_hd__conb_1
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_527_ net202 _101_ vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__ebufn_8
XFILLER_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_243_ net14 net21 net10 _046_ vssd1 vssd1 vccd1 vccd1 _047_ sky130_fd_sc_hd__a31o_1
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput18 io_in[34] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_2
X_174_ _091_ vssd1 vssd1 vccd1 vccd1 _110_ sky130_fd_sc_hd__inv_2
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_117 vssd1 vssd1 vccd1 vccd1 macro_decap_3_117/HI la_data_out[84] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_106 vssd1 vssd1 vccd1 vccd1 macro_decap_3_106/HI la_data_out[73] sky130_fd_sc_hd__conb_1
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_128 vssd1 vssd1 vccd1 vccd1 macro_decap_3_128/HI la_data_out[95] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_139 vssd1 vssd1 vccd1 vccd1 macro_decap_3_139/HI la_data_out[106] sky130_fd_sc_hd__conb_1
XFILLER_36_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_226_ net13 _022_ vssd1 vssd1 vccd1 vccd1 _033_ sky130_fd_sc_hd__and2_1
XFILLER_8_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_157_ net1 vssd1 vssd1 vccd1 vccd1 _124_ sky130_fd_sc_hd__inv_2
XFILLER_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__239__A2 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_209_ net9 _000_ _001_ vssd1 vssd1 vccd1 vccd1 _016_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__246__A _089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_524__199 vssd1 vssd1 vccd1 vccd1 _524__199/HI net199 sky130_fd_sc_hd__conb_1
XFILLER_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_543_ net218 _117_ vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__ebufn_8
XFILLER_17_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__211__B1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_190_ _092_ vssd1 vssd1 vccd1 vccd1 _095_ sky130_fd_sc_hd__inv_2
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_80 vssd1 vssd1 vccd1 vccd1 macro_decap_3_80/HI la_data_out[15] sky130_fd_sc_hd__conb_1
XFILLER_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_91 vssd1 vssd1 vccd1 vccd1 macro_decap_3_91/HI la_data_out[26] sky130_fd_sc_hd__conb_1
XFILLER_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_526_ net201 _100_ vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__ebufn_8
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_242_ net14 net10 _045_ vssd1 vssd1 vccd1 vccd1 _046_ sky130_fd_sc_hd__o21a_1
Xinput19 io_in[35] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_173_ _091_ vssd1 vssd1 vccd1 vccd1 _111_ sky130_fd_sc_hd__inv_2
XFILLER_10_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_107 vssd1 vssd1 vccd1 vccd1 macro_decap_3_107/HI la_data_out[74] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_118 vssd1 vssd1 vccd1 vccd1 macro_decap_3_118/HI la_data_out[85] sky130_fd_sc_hd__conb_1
XFILLER_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_129 vssd1 vssd1 vccd1 vccd1 macro_decap_3_129/HI la_data_out[96] sky130_fd_sc_hd__conb_1
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_225_ _029_ _030_ _031_ vssd1 vssd1 vccd1 vccd1 _032_ sky130_fd_sc_hd__a21o_1
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__159__A _089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_545__220 vssd1 vssd1 vccd1 vccd1 _545__220/HI net220 sky130_fd_sc_hd__conb_1
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_208_ _006_ _012_ _013_ _014_ vssd1 vssd1 vccd1 vccd1 _015_ sky130_fd_sc_hd__a211o_1
XFILLER_11_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_529__204 vssd1 vssd1 vccd1 vccd1 _529__204/HI net204 sky130_fd_sc_hd__conb_1
XFILLER_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_542_ net217 _116_ vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__ebufn_8
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_70 vssd1 vssd1 vccd1 vccd1 macro_decap_3_70/HI la_data_out[5] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_81 vssd1 vssd1 vccd1 vccd1 macro_decap_3_81/HI la_data_out[16] sky130_fd_sc_hd__conb_1
XFILLER_92_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_92 vssd1 vssd1 vccd1 vccd1 macro_decap_3_92/HI la_data_out[27] sky130_fd_sc_hd__conb_1
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_525_ net200 _099_ vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__ebufn_8
XFILLER_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__269__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_241_ net14 net10 _044_ net20 vssd1 vssd1 vccd1 vccd1 _045_ sky130_fd_sc_hd__o2bb2a_1
X_172_ _091_ vssd1 vssd1 vccd1 vccd1 _112_ sky130_fd_sc_hd__inv_2
XFILLER_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_108 vssd1 vssd1 vccd1 vccd1 macro_decap_3_108/HI la_data_out[75] sky130_fd_sc_hd__conb_1
XFILLER_56_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_119 vssd1 vssd1 vccd1 vccd1 macro_decap_3_119/HI la_data_out[86] sky130_fd_sc_hd__conb_1
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__265__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_224_ net11 _027_ _028_ vssd1 vssd1 vccd1 vccd1 _031_ sky130_fd_sc_hd__and3_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_207_ net4 _005_ vssd1 vssd1 vccd1 vccd1 _014_ sky130_fd_sc_hd__and2_1
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_541_ net216 _115_ vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__ebufn_8
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_60 vssd1 vssd1 vccd1 vccd1 macro_decap_3_60/HI io_out[33] sky130_fd_sc_hd__conb_1
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_71 vssd1 vssd1 vccd1 vccd1 macro_decap_3_71/HI la_data_out[6] sky130_fd_sc_hd__conb_1
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_82 vssd1 vssd1 vccd1 vccd1 macro_decap_3_82/HI la_data_out[17] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_93 vssd1 vssd1 vccd1 vccd1 macro_decap_3_93/HI la_data_out[28] sky130_fd_sc_hd__conb_1
XANTENNA_input11_A io_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_524_ net199 _098_ vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__ebufn_8
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input3_A io_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_240_ net21 vssd1 vssd1 vccd1 vccd1 _044_ sky130_fd_sc_hd__inv_2
XFILLER_52_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_171_ _091_ vssd1 vssd1 vccd1 vccd1 _113_ sky130_fd_sc_hd__inv_2
XFILLER_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_109 vssd1 vssd1 vccd1 vccd1 macro_decap_3_109/HI la_data_out[76] sky130_fd_sc_hd__conb_1
XFILLER_83_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_223_ net10 net14 vssd1 vssd1 vccd1 vccd1 _030_ sky130_fd_sc_hd__or2b_1
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__276__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_206_ net5 _002_ vssd1 vssd1 vccd1 vccd1 _013_ sky130_fd_sc_hd__and2_1
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_535__210 vssd1 vssd1 vccd1 vccd1 _535__210/HI net210 sky130_fd_sc_hd__conb_1
XFILLER_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_540_ net215 _114_ vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__ebufn_8
XFILLER_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xmacro_decap_3_61 vssd1 vssd1 vccd1 vccd1 macro_decap_3_61/HI io_out[34] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_50 vssd1 vssd1 vccd1 vccd1 macro_decap_3_50/HI io_out[23] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_72 vssd1 vssd1 vccd1 vccd1 macro_decap_3_72/HI la_data_out[7] sky130_fd_sc_hd__conb_1
XFILLER_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xmacro_decap_3_83 vssd1 vssd1 vccd1 vccd1 macro_decap_3_83/HI la_data_out[18] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_94 vssd1 vssd1 vccd1 vccd1 macro_decap_3_94/HI la_data_out[29] sky130_fd_sc_hd__conb_1
XFILLER_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_523_ net198 _097_ vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__ebufn_8
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__284__A net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_170_ _089_ vssd1 vssd1 vccd1 vccd1 _091_ sky130_fd_sc_hd__buf_4
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_222_ _027_ _028_ net11 vssd1 vssd1 vccd1 vccd1 _029_ sky130_fd_sc_hd__a21o_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_205_ _009_ _010_ _011_ vssd1 vssd1 vccd1 vccd1 _012_ sky130_fd_sc_hd__a21o_1
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_40 vssd1 vssd1 vccd1 vccd1 macro_decap_3_40/HI io_oeb[36] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_62 vssd1 vssd1 vccd1 vccd1 macro_decap_3_62/HI io_out[35] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_51 vssd1 vssd1 vccd1 vccd1 macro_decap_3_51/HI io_out[24] sky130_fd_sc_hd__conb_1
XFILLER_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_73 vssd1 vssd1 vccd1 vccd1 macro_decap_3_73/HI la_data_out[8] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_84 vssd1 vssd1 vccd1 vccd1 macro_decap_3_84/HI la_data_out[19] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_95 vssd1 vssd1 vccd1 vccd1 macro_decap_3_95/HI la_data_out[30] sky130_fd_sc_hd__conb_1
XFILLER_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_522_ net197 _096_ vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__ebufn_8
XFILLER_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_520__195 vssd1 vssd1 vccd1 vccd1 _520__195/HI net195 sky130_fd_sc_hd__conb_1
XFILLER_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_221_ net14 _020_ net15 vssd1 vssd1 vccd1 vccd1 _028_ sky130_fd_sc_hd__a21bo_1
XFILLER_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_204_ net3 _007_ _008_ vssd1 vssd1 vccd1 vccd1 _011_ sky130_fd_sc_hd__and3_1
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_250 vssd1 vssd1 vccd1 vccd1 macro_decap_3_250/HI io_oeb[24] sky130_fd_sc_hd__conb_1
XFILLER_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_41 vssd1 vssd1 vccd1 vccd1 macro_decap_3_41/HI io_oeb[37] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_63 vssd1 vssd1 vccd1 vccd1 macro_decap_3_63/HI io_out[36] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_52 vssd1 vssd1 vccd1 vccd1 macro_decap_3_52/HI io_out[25] sky130_fd_sc_hd__conb_1
XFILLER_92_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_74 vssd1 vssd1 vccd1 vccd1 macro_decap_3_74/HI la_data_out[9] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_85 vssd1 vssd1 vccd1 vccd1 macro_decap_3_85/HI la_data_out[20] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_96 vssd1 vssd1 vccd1 vccd1 macro_decap_3_96/HI la_data_out[31] sky130_fd_sc_hd__conb_1
XFILLER_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_521_ net196 _095_ vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__ebufn_8
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_525__200 vssd1 vssd1 vccd1 vccd1 _525__200/HI net200 sky130_fd_sc_hd__conb_1
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input1_A io_active vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_220_ net15 _020_ net14 vssd1 vssd1 vccd1 vccd1 _027_ sky130_fd_sc_hd__nand3b_1
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_203_ net2 net6 vssd1 vssd1 vccd1 vccd1 _010_ sky130_fd_sc_hd__or2b_1
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__235__B1 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmacro_decap_3_240 vssd1 vssd1 vccd1 vccd1 macro_decap_3_240/HI io_oeb[14] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_251 vssd1 vssd1 vccd1 vccd1 macro_decap_3_251/HI io_oeb[25] sky130_fd_sc_hd__conb_1
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_542__217 vssd1 vssd1 vccd1 vccd1 _542__217/HI net217 sky130_fd_sc_hd__conb_1
XFILLER_25_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_53 vssd1 vssd1 vccd1 vccd1 macro_decap_3_53/HI io_out[26] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_42 vssd1 vssd1 vccd1 vccd1 macro_decap_3_42/HI io_out[1] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_64 vssd1 vssd1 vccd1 vccd1 macro_decap_3_64/HI io_out[37] sky130_fd_sc_hd__conb_1
XFILLER_66_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmacro_decap_3_86 vssd1 vssd1 vccd1 vccd1 macro_decap_3_86/HI la_data_out[21] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_75 vssd1 vssd1 vccd1 vccd1 macro_decap_3_75/HI la_data_out[10] sky130_fd_sc_hd__conb_1
X_520_ net195 _094_ vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__ebufn_8
Xmacro_decap_3_97 vssd1 vssd1 vccd1 vccd1 macro_decap_3_97/HI la_data_out[64] sky130_fd_sc_hd__conb_1
XFILLER_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_548__223 vssd1 vssd1 vccd1 vccd1 _548__223/HI net223 sky130_fd_sc_hd__conb_1
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_296_ _079_ _082_ _088_ net26 net30 vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__o32a_1
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_279_ _075_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__253__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_202_ _007_ _008_ net3 vssd1 vssd1 vccd1 vccd1 _009_ sky130_fd_sc_hd__a21o_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_230 vssd1 vssd1 vccd1 vccd1 macro_decap_3_230/HI io_oeb[4] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_241 vssd1 vssd1 vccd1 vccd1 macro_decap_3_241/HI io_oeb[15] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_252 vssd1 vssd1 vccd1 vccd1 macro_decap_3_252/HI io_oeb[26] sky130_fd_sc_hd__conb_1
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xmacro_decap_3_43 vssd1 vssd1 vccd1 vccd1 macro_decap_3_43/HI io_out[2] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_54 vssd1 vssd1 vccd1 vccd1 macro_decap_3_54/HI io_out[27] sky130_fd_sc_hd__conb_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmacro_decap_3_76 vssd1 vssd1 vccd1 vccd1 macro_decap_3_76/HI la_data_out[11] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_65 vssd1 vssd1 vccd1 vccd1 macro_decap_3_65/HI la_data_out[0] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_87 vssd1 vssd1 vccd1 vccd1 macro_decap_3_87/HI la_data_out[22] sky130_fd_sc_hd__conb_1
XFILLER_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_98 vssd1 vssd1 vccd1 vccd1 macro_decap_3_98/HI la_data_out[65] sky130_fd_sc_hd__conb_1
XFILLER_57_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_295_ net19 _078_ _080_ _081_ _089_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__o221a_1
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_278_ _089_ _067_ vssd1 vssd1 vccd1 vccd1 _075_ sky130_fd_sc_hd__and2_1
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_68_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_201_ net6 _000_ net7 vssd1 vssd1 vccd1 vccd1 _008_ sky130_fd_sc_hd__a21bo_1
XFILLER_90_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_253 vssd1 vssd1 vccd1 vccd1 macro_decap_3_253/HI io_oeb[27] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_231 vssd1 vssd1 vccd1 vccd1 macro_decap_3_231/HI io_oeb[5] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_242 vssd1 vssd1 vccd1 vccd1 macro_decap_3_242/HI io_oeb[16] sky130_fd_sc_hd__conb_1
XFILLER_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_44 vssd1 vssd1 vccd1 vccd1 macro_decap_3_44/HI io_out[3] sky130_fd_sc_hd__conb_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmacro_decap_3_55 vssd1 vssd1 vccd1 vccd1 macro_decap_3_55/HI io_out[28] sky130_fd_sc_hd__conb_1
XFILLER_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmacro_decap_3_66 vssd1 vssd1 vccd1 vccd1 macro_decap_3_66/HI la_data_out[1] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_77 vssd1 vssd1 vccd1 vccd1 macro_decap_3_77/HI la_data_out[12] sky130_fd_sc_hd__conb_1
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xmacro_decap_3_88 vssd1 vssd1 vccd1 vccd1 macro_decap_3_88/HI la_data_out[23] sky130_fd_sc_hd__conb_1
Xmacro_decap_3_99 vssd1 vssd1 vccd1 vccd1 macro_decap_3_99/HI la_data_out[66] sky130_fd_sc_hd__conb_1
XFILLER_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_2
XFILLER_95_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_532__207 vssd1 vssd1 vccd1 vccd1 _532__207/HI net207 sky130_fd_sc_hd__conb_1
XFILLER_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
.ends

