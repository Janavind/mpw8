// This is the unpowered netlist.
module macro_7 (io_active,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input io_active;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net228;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net229;
 wire net257;
 wire net258;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net46;
 wire net47;
 wire net43;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net44;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net45;
 wire net66;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net76;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net77;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net67;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net68;
 wire net96;
 wire net97;
 wire net69;
 wire net70;
 wire net71;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net72;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net73;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net74;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net75;
 wire net162;
 wire net163;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net164;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net165;
 wire net193;
 wire net194;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;

 sky130_fd_sc_hd__clkinv_2 _157_ (.A(net1),
    .Y(_124_));
 sky130_fd_sc_hd__buf_4 _158_ (.A(net1),
    .X(_089_));
 sky130_fd_sc_hd__buf_4 _159_ (.A(_089_),
    .X(_090_));
 sky130_fd_sc_hd__inv_2 _160_ (.A(_090_),
    .Y(_123_));
 sky130_fd_sc_hd__inv_2 _161_ (.A(_090_),
    .Y(_122_));
 sky130_fd_sc_hd__inv_2 _162_ (.A(_090_),
    .Y(_121_));
 sky130_fd_sc_hd__inv_2 _163_ (.A(_090_),
    .Y(_120_));
 sky130_fd_sc_hd__inv_2 _164_ (.A(_090_),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _165_ (.A(_090_),
    .Y(_118_));
 sky130_fd_sc_hd__inv_2 _166_ (.A(_090_),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _167_ (.A(_090_),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _168_ (.A(_090_),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _169_ (.A(_090_),
    .Y(_114_));
 sky130_fd_sc_hd__buf_4 _170_ (.A(_089_),
    .X(_091_));
 sky130_fd_sc_hd__inv_2 _171_ (.A(_091_),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _172_ (.A(_091_),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _173_ (.A(_091_),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _174_ (.A(_091_),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _175_ (.A(_091_),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _176_ (.A(_091_),
    .Y(_108_));
 sky130_fd_sc_hd__inv_2 _177_ (.A(_091_),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _178_ (.A(_091_),
    .Y(_106_));
 sky130_fd_sc_hd__inv_2 _179_ (.A(_091_),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _180_ (.A(_091_),
    .Y(_104_));
 sky130_fd_sc_hd__buf_4 _181_ (.A(_089_),
    .X(_092_));
 sky130_fd_sc_hd__inv_2 _182_ (.A(_092_),
    .Y(_103_));
 sky130_fd_sc_hd__inv_2 _183_ (.A(_092_),
    .Y(_102_));
 sky130_fd_sc_hd__inv_2 _184_ (.A(_092_),
    .Y(_101_));
 sky130_fd_sc_hd__inv_2 _185_ (.A(_092_),
    .Y(_100_));
 sky130_fd_sc_hd__inv_2 _186_ (.A(_092_),
    .Y(_099_));
 sky130_fd_sc_hd__inv_2 _187_ (.A(_092_),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _188_ (.A(_092_),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _189_ (.A(_092_),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _190_ (.A(_092_),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _191_ (.A(_092_),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _192_ (.A(_089_),
    .Y(_093_));
 sky130_fd_sc_hd__nand2b_1 _193_ (.A_N(net19),
    .B(net18),
    .Y(_000_));
 sky130_fd_sc_hd__o31a_1 _194_ (.A1(net8),
    .A2(net6),
    .A3(net7),
    .B1(_000_),
    .X(_001_));
 sky130_fd_sc_hd__xnor2_1 _195_ (.A(net9),
    .B(_001_),
    .Y(_002_));
 sky130_fd_sc_hd__or2_1 _196_ (.A(net5),
    .B(_002_),
    .X(_003_));
 sky130_fd_sc_hd__o21a_1 _197_ (.A1(net6),
    .A2(net7),
    .B1(_000_),
    .X(_004_));
 sky130_fd_sc_hd__xnor2_1 _198_ (.A(net8),
    .B(_004_),
    .Y(_005_));
 sky130_fd_sc_hd__or2_1 _199_ (.A(net4),
    .B(_005_),
    .X(_006_));
 sky130_fd_sc_hd__nand3b_1 _200_ (.A_N(net7),
    .B(_000_),
    .C(net6),
    .Y(_007_));
 sky130_fd_sc_hd__a21bo_1 _201_ (.A1(net6),
    .A2(_000_),
    .B1_N(net7),
    .X(_008_));
 sky130_fd_sc_hd__a21o_1 _202_ (.A1(_007_),
    .A2(_008_),
    .B1(net3),
    .X(_009_));
 sky130_fd_sc_hd__or2b_1 _203_ (.A(net2),
    .B_N(net6),
    .X(_010_));
 sky130_fd_sc_hd__and3_1 _204_ (.A(net3),
    .B(_007_),
    .C(_008_),
    .X(_011_));
 sky130_fd_sc_hd__a21o_1 _205_ (.A1(_009_),
    .A2(_010_),
    .B1(_011_),
    .X(_012_));
 sky130_fd_sc_hd__and2_1 _206_ (.A(net5),
    .B(_002_),
    .X(_013_));
 sky130_fd_sc_hd__and2_1 _207_ (.A(net4),
    .B(_005_),
    .X(_014_));
 sky130_fd_sc_hd__a211o_1 _208_ (.A1(_006_),
    .A2(_012_),
    .B1(_013_),
    .C1(_014_),
    .X(_015_));
 sky130_fd_sc_hd__a21oi_1 _209_ (.A1(net9),
    .A2(_000_),
    .B1(_001_),
    .Y(_016_));
 sky130_fd_sc_hd__a21oi_1 _210_ (.A1(_003_),
    .A2(_015_),
    .B1(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__a31o_1 _211_ (.A1(_016_),
    .A2(_003_),
    .A3(_015_),
    .B1(net19),
    .X(_018_));
 sky130_fd_sc_hd__or2_1 _212_ (.A(_017_),
    .B(_018_),
    .X(_019_));
 sky130_fd_sc_hd__nand2b_1 _213_ (.A_N(net21),
    .B(net20),
    .Y(_020_));
 sky130_fd_sc_hd__o31a_1 _214_ (.A1(net16),
    .A2(net14),
    .A3(net15),
    .B1(_020_),
    .X(_021_));
 sky130_fd_sc_hd__xnor2_1 _215_ (.A(net17),
    .B(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__or2_1 _216_ (.A(net13),
    .B(_022_),
    .X(_023_));
 sky130_fd_sc_hd__o21a_1 _217_ (.A1(net14),
    .A2(net15),
    .B1(_020_),
    .X(_024_));
 sky130_fd_sc_hd__xnor2_1 _218_ (.A(net16),
    .B(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__or2_1 _219_ (.A(net12),
    .B(_025_),
    .X(_026_));
 sky130_fd_sc_hd__nand3b_1 _220_ (.A_N(net15),
    .B(_020_),
    .C(net14),
    .Y(_027_));
 sky130_fd_sc_hd__a21bo_1 _221_ (.A1(net14),
    .A2(_020_),
    .B1_N(net15),
    .X(_028_));
 sky130_fd_sc_hd__a21o_1 _222_ (.A1(_027_),
    .A2(_028_),
    .B1(net11),
    .X(_029_));
 sky130_fd_sc_hd__or2b_1 _223_ (.A(net10),
    .B_N(net14),
    .X(_030_));
 sky130_fd_sc_hd__and3_1 _224_ (.A(net11),
    .B(_027_),
    .C(_028_),
    .X(_031_));
 sky130_fd_sc_hd__a21o_1 _225_ (.A1(_029_),
    .A2(_030_),
    .B1(_031_),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _226_ (.A(net13),
    .B(_022_),
    .X(_033_));
 sky130_fd_sc_hd__and2_1 _227_ (.A(net12),
    .B(_025_),
    .X(_034_));
 sky130_fd_sc_hd__a211o_1 _228_ (.A1(_026_),
    .A2(_032_),
    .B1(_033_),
    .C1(_034_),
    .X(_035_));
 sky130_fd_sc_hd__a21oi_1 _229_ (.A1(net17),
    .A2(_020_),
    .B1(_021_),
    .Y(_036_));
 sky130_fd_sc_hd__a21oi_1 _230_ (.A1(_023_),
    .A2(_035_),
    .B1(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__a31o_1 _231_ (.A1(_036_),
    .A2(_023_),
    .A3(_035_),
    .B1(net21),
    .X(_038_));
 sky130_fd_sc_hd__or2_1 _232_ (.A(_037_),
    .B(_038_),
    .X(_039_));
 sky130_fd_sc_hd__nor3_2 _233_ (.A(_124_),
    .B(_037_),
    .C(_038_),
    .Y(net31));
 sky130_fd_sc_hd__nor3_1 _234_ (.A(_124_),
    .B(_017_),
    .C(_018_),
    .Y(net32));
 sky130_fd_sc_hd__o22a_1 _235_ (.A1(_019_),
    .A2(_039_),
    .B1(net31),
    .B2(net32),
    .X(net22));
 sky130_fd_sc_hd__inv_2 _236_ (.A(net19),
    .Y(_040_));
 sky130_fd_sc_hd__o2bb2a_1 _237_ (.A1_N(net6),
    .A2_N(net2),
    .B1(_040_),
    .B2(net18),
    .X(_041_));
 sky130_fd_sc_hd__o21a_1 _238_ (.A1(net6),
    .A2(net2),
    .B1(_041_),
    .X(_042_));
 sky130_fd_sc_hd__a31o_1 _239_ (.A1(net6),
    .A2(net19),
    .A3(net2),
    .B1(_042_),
    .X(_043_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(net21),
    .Y(_044_));
 sky130_fd_sc_hd__o2bb2a_1 _241_ (.A1_N(net14),
    .A2_N(net10),
    .B1(_044_),
    .B2(net20),
    .X(_045_));
 sky130_fd_sc_hd__o21a_1 _242_ (.A1(net14),
    .A2(net10),
    .B1(_045_),
    .X(_046_));
 sky130_fd_sc_hd__a31o_1 _243_ (.A1(net14),
    .A2(net21),
    .A3(net10),
    .B1(_046_),
    .X(_047_));
 sky130_fd_sc_hd__and2_1 _244_ (.A(_089_),
    .B(_047_),
    .X(_048_));
 sky130_fd_sc_hd__clkbuf_1 _245_ (.A(_048_),
    .X(net23));
 sky130_fd_sc_hd__and2_1 _246_ (.A(_089_),
    .B(_043_),
    .X(_049_));
 sky130_fd_sc_hd__clkbuf_1 _247_ (.A(_049_),
    .X(net27));
 sky130_fd_sc_hd__o2bb2a_1 _248_ (.A1_N(_043_),
    .A2_N(_047_),
    .B1(net23),
    .B2(net27),
    .X(net33));
 sky130_fd_sc_hd__or2b_1 _249_ (.A(_011_),
    .B_N(_009_),
    .X(_050_));
 sky130_fd_sc_hd__xnor2_1 _250_ (.A(_050_),
    .B(_010_),
    .Y(_051_));
 sky130_fd_sc_hd__o21a_1 _251_ (.A1(net7),
    .A2(net18),
    .B1(net3),
    .X(_052_));
 sky130_fd_sc_hd__a211o_1 _252_ (.A1(net7),
    .A2(net18),
    .B1(_040_),
    .C1(_052_),
    .X(_053_));
 sky130_fd_sc_hd__o21a_1 _253_ (.A1(net19),
    .A2(_051_),
    .B1(_053_),
    .X(_054_));
 sky130_fd_sc_hd__or2b_1 _254_ (.A(_031_),
    .B_N(_029_),
    .X(_055_));
 sky130_fd_sc_hd__xnor2_1 _255_ (.A(_055_),
    .B(_030_),
    .Y(_056_));
 sky130_fd_sc_hd__o21a_1 _256_ (.A1(net15),
    .A2(net20),
    .B1(net11),
    .X(_057_));
 sky130_fd_sc_hd__a211o_1 _257_ (.A1(net15),
    .A2(net20),
    .B1(_044_),
    .C1(_057_),
    .X(_058_));
 sky130_fd_sc_hd__o21a_1 _258_ (.A1(net21),
    .A2(_056_),
    .B1(_058_),
    .X(_059_));
 sky130_fd_sc_hd__and2_1 _259_ (.A(_089_),
    .B(_059_),
    .X(_060_));
 sky130_fd_sc_hd__clkbuf_1 _260_ (.A(_060_),
    .X(net24));
 sky130_fd_sc_hd__and2_1 _261_ (.A(_089_),
    .B(_054_),
    .X(_061_));
 sky130_fd_sc_hd__clkbuf_1 _262_ (.A(_061_),
    .X(net28));
 sky130_fd_sc_hd__o2bb2a_1 _263_ (.A1_N(_054_),
    .A2_N(_059_),
    .B1(net24),
    .B2(net28),
    .X(net34));
 sky130_fd_sc_hd__a21o_1 _264_ (.A1(net18),
    .A2(net4),
    .B1(net8),
    .X(_062_));
 sky130_fd_sc_hd__or2_1 _265_ (.A(net18),
    .B(net4),
    .X(_063_));
 sky130_fd_sc_hd__xor2_1 _266_ (.A(net4),
    .B(_005_),
    .X(_064_));
 sky130_fd_sc_hd__or2_1 _267_ (.A(_064_),
    .B(_012_),
    .X(_065_));
 sky130_fd_sc_hd__a21oi_1 _268_ (.A1(_064_),
    .A2(_012_),
    .B1(net19),
    .Y(_066_));
 sky130_fd_sc_hd__a32o_1 _269_ (.A1(net19),
    .A2(_062_),
    .A3(_063_),
    .B1(_065_),
    .B2(_066_),
    .X(_067_));
 sky130_fd_sc_hd__a21o_1 _270_ (.A1(net20),
    .A2(net12),
    .B1(net16),
    .X(_068_));
 sky130_fd_sc_hd__or2_1 _271_ (.A(net20),
    .B(net12),
    .X(_069_));
 sky130_fd_sc_hd__xor2_1 _272_ (.A(net12),
    .B(_025_),
    .X(_070_));
 sky130_fd_sc_hd__or2_1 _273_ (.A(_070_),
    .B(_032_),
    .X(_071_));
 sky130_fd_sc_hd__a21oi_1 _274_ (.A1(_070_),
    .A2(_032_),
    .B1(net21),
    .Y(_072_));
 sky130_fd_sc_hd__a32o_1 _275_ (.A1(net21),
    .A2(_068_),
    .A3(_069_),
    .B1(_071_),
    .B2(_072_),
    .X(_073_));
 sky130_fd_sc_hd__and2_1 _276_ (.A(net1),
    .B(_073_),
    .X(_074_));
 sky130_fd_sc_hd__clkbuf_1 _277_ (.A(_074_),
    .X(net25));
 sky130_fd_sc_hd__and2_1 _278_ (.A(_089_),
    .B(_067_),
    .X(_075_));
 sky130_fd_sc_hd__clkbuf_1 _279_ (.A(_075_),
    .X(net29));
 sky130_fd_sc_hd__o2bb2a_1 _280_ (.A1_N(_067_),
    .A2_N(_073_),
    .B1(net25),
    .B2(net29),
    .X(net35));
 sky130_fd_sc_hd__a21oi_1 _281_ (.A1(_006_),
    .A2(_012_),
    .B1(_014_),
    .Y(_076_));
 sky130_fd_sc_hd__and2b_1 _282_ (.A_N(_013_),
    .B(_003_),
    .X(_077_));
 sky130_fd_sc_hd__xnor2_1 _283_ (.A(_076_),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__nor2_1 _284_ (.A(net19),
    .B(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__o21a_1 _285_ (.A1(net9),
    .A2(net18),
    .B1(net5),
    .X(_080_));
 sky130_fd_sc_hd__a21o_1 _286_ (.A1(net9),
    .A2(net18),
    .B1(_040_),
    .X(_081_));
 sky130_fd_sc_hd__nor2_1 _287_ (.A(_080_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__a21o_1 _288_ (.A1(_026_),
    .A2(_032_),
    .B1(_034_),
    .X(_083_));
 sky130_fd_sc_hd__and2b_1 _289_ (.A_N(_033_),
    .B(_023_),
    .X(_084_));
 sky130_fd_sc_hd__xnor2_1 _290_ (.A(_083_),
    .B(_084_),
    .Y(_085_));
 sky130_fd_sc_hd__o21a_1 _291_ (.A1(net17),
    .A2(net20),
    .B1(net13),
    .X(_086_));
 sky130_fd_sc_hd__a211oi_2 _292_ (.A1(net17),
    .A2(net20),
    .B1(_044_),
    .C1(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__a21o_1 _293_ (.A1(_044_),
    .A2(_085_),
    .B1(_087_),
    .X(_088_));
 sky130_fd_sc_hd__a211oi_2 _294_ (.A1(_044_),
    .A2(_085_),
    .B1(_087_),
    .C1(_124_),
    .Y(net26));
 sky130_fd_sc_hd__o221a_1 _295_ (.A1(net19),
    .A2(_078_),
    .B1(_080_),
    .B2(_081_),
    .C1(_089_),
    .X(net30));
 sky130_fd_sc_hd__o32a_1 _296_ (.A1(_079_),
    .A2(_082_),
    .A3(_088_),
    .B1(net26),
    .B2(net30),
    .X(net36));
 sky130_fd_sc_hd__conb_1 macro_7_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 macro_7_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 macro_7_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 macro_7_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 macro_7_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 macro_7_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 macro_7_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 macro_7_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 macro_7_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 macro_7_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 macro_7_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 macro_7_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 macro_7_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 macro_7_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 macro_7_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 macro_7_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 macro_7_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 macro_7_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 macro_7_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 macro_7_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 macro_7_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 macro_7_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 macro_7_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 macro_7_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 macro_7_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 macro_7_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 macro_7_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 macro_7_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 macro_7_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 macro_7_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 macro_7_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 macro_7_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 macro_7_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 macro_7_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 macro_7_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 macro_7_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 macro_7_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 macro_7_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 macro_7_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 macro_7_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 macro_7_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 macro_7_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 macro_7_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 macro_7_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 macro_7_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 macro_7_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 macro_7_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 macro_7_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 macro_7_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 macro_7_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 macro_7_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 macro_7_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 macro_7_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 macro_7_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 macro_7_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 macro_7_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 macro_7_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 macro_7_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 macro_7_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 macro_7_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 macro_7_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 macro_7_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 macro_7_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 macro_7_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 macro_7_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 macro_7_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 macro_7_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 macro_7_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 macro_7_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 macro_7_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 macro_7_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 macro_7_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 macro_7_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 macro_7_111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 macro_7_112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 macro_7_113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 macro_7_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 macro_7_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 macro_7_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 macro_7_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 macro_7_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 macro_7_119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 macro_7_120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 macro_7_121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 macro_7_122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 macro_7_123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 macro_7_124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 macro_7_125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 macro_7_126 (.LO(net126));
 sky130_fd_sc_hd__conb_1 macro_7_127 (.LO(net127));
 sky130_fd_sc_hd__conb_1 macro_7_128 (.LO(net128));
 sky130_fd_sc_hd__conb_1 macro_7_129 (.LO(net129));
 sky130_fd_sc_hd__conb_1 macro_7_130 (.LO(net130));
 sky130_fd_sc_hd__conb_1 macro_7_131 (.LO(net131));
 sky130_fd_sc_hd__conb_1 macro_7_132 (.LO(net132));
 sky130_fd_sc_hd__conb_1 macro_7_133 (.LO(net133));
 sky130_fd_sc_hd__conb_1 macro_7_134 (.LO(net134));
 sky130_fd_sc_hd__conb_1 macro_7_135 (.LO(net135));
 sky130_fd_sc_hd__conb_1 macro_7_136 (.LO(net136));
 sky130_fd_sc_hd__conb_1 macro_7_137 (.LO(net137));
 sky130_fd_sc_hd__conb_1 macro_7_138 (.LO(net138));
 sky130_fd_sc_hd__conb_1 macro_7_139 (.LO(net139));
 sky130_fd_sc_hd__conb_1 macro_7_140 (.LO(net140));
 sky130_fd_sc_hd__conb_1 macro_7_141 (.LO(net141));
 sky130_fd_sc_hd__conb_1 macro_7_142 (.LO(net142));
 sky130_fd_sc_hd__conb_1 macro_7_143 (.LO(net143));
 sky130_fd_sc_hd__conb_1 macro_7_144 (.LO(net144));
 sky130_fd_sc_hd__conb_1 macro_7_145 (.LO(net145));
 sky130_fd_sc_hd__conb_1 macro_7_146 (.LO(net146));
 sky130_fd_sc_hd__conb_1 macro_7_147 (.LO(net147));
 sky130_fd_sc_hd__conb_1 macro_7_148 (.LO(net148));
 sky130_fd_sc_hd__conb_1 macro_7_149 (.LO(net149));
 sky130_fd_sc_hd__conb_1 macro_7_150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 macro_7_151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 macro_7_152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 macro_7_153 (.LO(net153));
 sky130_fd_sc_hd__conb_1 macro_7_154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 macro_7_155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 macro_7_156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 macro_7_157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 macro_7_158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 macro_7_159 (.LO(net159));
 sky130_fd_sc_hd__conb_1 macro_7_160 (.LO(net160));
 sky130_fd_sc_hd__conb_1 macro_7_161 (.LO(net161));
 sky130_fd_sc_hd__conb_1 macro_7_162 (.LO(net162));
 sky130_fd_sc_hd__conb_1 macro_7_163 (.LO(net163));
 sky130_fd_sc_hd__conb_1 macro_7_164 (.LO(net164));
 sky130_fd_sc_hd__conb_1 macro_7_165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 macro_7_166 (.LO(net166));
 sky130_fd_sc_hd__conb_1 macro_7_167 (.LO(net167));
 sky130_fd_sc_hd__conb_1 macro_7_168 (.LO(net168));
 sky130_fd_sc_hd__conb_1 macro_7_169 (.LO(net169));
 sky130_fd_sc_hd__conb_1 macro_7_170 (.LO(net170));
 sky130_fd_sc_hd__conb_1 macro_7_171 (.LO(net171));
 sky130_fd_sc_hd__conb_1 macro_7_172 (.LO(net172));
 sky130_fd_sc_hd__conb_1 macro_7_173 (.LO(net173));
 sky130_fd_sc_hd__conb_1 macro_7_174 (.LO(net174));
 sky130_fd_sc_hd__conb_1 macro_7_175 (.LO(net175));
 sky130_fd_sc_hd__conb_1 macro_7_176 (.LO(net176));
 sky130_fd_sc_hd__conb_1 macro_7_177 (.LO(net177));
 sky130_fd_sc_hd__conb_1 macro_7_178 (.LO(net178));
 sky130_fd_sc_hd__conb_1 macro_7_179 (.LO(net179));
 sky130_fd_sc_hd__conb_1 macro_7_180 (.LO(net180));
 sky130_fd_sc_hd__conb_1 macro_7_181 (.LO(net181));
 sky130_fd_sc_hd__conb_1 macro_7_182 (.LO(net182));
 sky130_fd_sc_hd__conb_1 macro_7_183 (.LO(net183));
 sky130_fd_sc_hd__conb_1 macro_7_184 (.LO(net184));
 sky130_fd_sc_hd__conb_1 macro_7_185 (.LO(net185));
 sky130_fd_sc_hd__conb_1 macro_7_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 macro_7_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 macro_7_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 macro_7_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 macro_7_190 (.LO(net190));
 sky130_fd_sc_hd__conb_1 macro_7_191 (.LO(net191));
 sky130_fd_sc_hd__conb_1 macro_7_192 (.LO(net192));
 sky130_fd_sc_hd__conb_1 macro_7_193 (.LO(net193));
 sky130_fd_sc_hd__conb_1 _519__194 (.LO(net194));
 sky130_fd_sc_hd__conb_1 _520__195 (.LO(net195));
 sky130_fd_sc_hd__conb_1 _521__196 (.LO(net196));
 sky130_fd_sc_hd__conb_1 _522__197 (.LO(net197));
 sky130_fd_sc_hd__conb_1 _523__198 (.LO(net198));
 sky130_fd_sc_hd__conb_1 _524__199 (.LO(net199));
 sky130_fd_sc_hd__conb_1 _525__200 (.LO(net200));
 sky130_fd_sc_hd__conb_1 _526__201 (.LO(net201));
 sky130_fd_sc_hd__conb_1 _527__202 (.LO(net202));
 sky130_fd_sc_hd__conb_1 _528__203 (.LO(net203));
 sky130_fd_sc_hd__conb_1 _529__204 (.LO(net204));
 sky130_fd_sc_hd__conb_1 _530__205 (.LO(net205));
 sky130_fd_sc_hd__conb_1 _531__206 (.LO(net206));
 sky130_fd_sc_hd__conb_1 _532__207 (.LO(net207));
 sky130_fd_sc_hd__conb_1 _533__208 (.LO(net208));
 sky130_fd_sc_hd__conb_1 _534__209 (.LO(net209));
 sky130_fd_sc_hd__conb_1 _535__210 (.LO(net210));
 sky130_fd_sc_hd__conb_1 _536__211 (.LO(net211));
 sky130_fd_sc_hd__conb_1 _537__212 (.LO(net212));
 sky130_fd_sc_hd__conb_1 _538__213 (.LO(net213));
 sky130_fd_sc_hd__conb_1 _539__214 (.LO(net214));
 sky130_fd_sc_hd__conb_1 _540__215 (.LO(net215));
 sky130_fd_sc_hd__conb_1 _541__216 (.LO(net216));
 sky130_fd_sc_hd__conb_1 _542__217 (.LO(net217));
 sky130_fd_sc_hd__conb_1 _543__218 (.LO(net218));
 sky130_fd_sc_hd__conb_1 _544__219 (.LO(net219));
 sky130_fd_sc_hd__conb_1 _545__220 (.LO(net220));
 sky130_fd_sc_hd__conb_1 _546__221 (.LO(net221));
 sky130_fd_sc_hd__conb_1 _547__222 (.LO(net222));
 sky130_fd_sc_hd__conb_1 _548__223 (.LO(net223));
 sky130_fd_sc_hd__conb_1 _549__224 (.LO(net224));
 sky130_fd_sc_hd__conb_1 _550__225 (.LO(net225));
 sky130_fd_sc_hd__conb_1 macro_7_226 (.LO(net226));
 sky130_fd_sc_hd__conb_1 macro_7_227 (.LO(net227));
 sky130_fd_sc_hd__conb_1 macro_7_228 (.LO(net228));
 sky130_fd_sc_hd__conb_1 macro_7_229 (.LO(net229));
 sky130_fd_sc_hd__conb_1 macro_7_230 (.LO(net230));
 sky130_fd_sc_hd__conb_1 macro_7_231 (.LO(net231));
 sky130_fd_sc_hd__conb_1 macro_7_232 (.LO(net232));
 sky130_fd_sc_hd__conb_1 macro_7_233 (.LO(net233));
 sky130_fd_sc_hd__conb_1 macro_7_234 (.LO(net234));
 sky130_fd_sc_hd__conb_1 macro_7_235 (.LO(net235));
 sky130_fd_sc_hd__conb_1 macro_7_236 (.LO(net236));
 sky130_fd_sc_hd__conb_1 macro_7_237 (.LO(net237));
 sky130_fd_sc_hd__conb_1 macro_7_238 (.LO(net238));
 sky130_fd_sc_hd__conb_1 macro_7_239 (.LO(net239));
 sky130_fd_sc_hd__conb_1 macro_7_240 (.LO(net240));
 sky130_fd_sc_hd__conb_1 macro_7_241 (.LO(net241));
 sky130_fd_sc_hd__conb_1 macro_7_242 (.LO(net242));
 sky130_fd_sc_hd__conb_1 macro_7_243 (.LO(net243));
 sky130_fd_sc_hd__conb_1 macro_7_244 (.LO(net244));
 sky130_fd_sc_hd__conb_1 macro_7_245 (.LO(net245));
 sky130_fd_sc_hd__conb_1 macro_7_246 (.LO(net246));
 sky130_fd_sc_hd__conb_1 macro_7_247 (.LO(net247));
 sky130_fd_sc_hd__conb_1 macro_7_248 (.LO(net248));
 sky130_fd_sc_hd__conb_1 macro_7_249 (.LO(net249));
 sky130_fd_sc_hd__conb_1 macro_7_250 (.LO(net250));
 sky130_fd_sc_hd__conb_1 macro_7_251 (.LO(net251));
 sky130_fd_sc_hd__conb_1 macro_7_252 (.LO(net252));
 sky130_fd_sc_hd__conb_1 macro_7_253 (.LO(net253));
 sky130_fd_sc_hd__conb_1 macro_7_254 (.LO(net254));
 sky130_fd_sc_hd__conb_1 macro_7_255 (.LO(net255));
 sky130_fd_sc_hd__conb_1 macro_7_256 (.LO(net256));
 sky130_fd_sc_hd__conb_1 macro_7_257 (.LO(net257));
 sky130_fd_sc_hd__conb_1 macro_7_258 (.LO(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__C1 (.DIODE(_089_));
 sky130_fd_sc_hd__ebufn_8 _519_ (.A(net194),
    .TE_B(_093_),
    .Z(la_data_out[32]));
 sky130_fd_sc_hd__ebufn_8 _520_ (.A(net195),
    .TE_B(_094_),
    .Z(la_data_out[33]));
 sky130_fd_sc_hd__ebufn_8 _521_ (.A(net196),
    .TE_B(_095_),
    .Z(la_data_out[34]));
 sky130_fd_sc_hd__ebufn_8 _522_ (.A(net197),
    .TE_B(_096_),
    .Z(la_data_out[35]));
 sky130_fd_sc_hd__ebufn_8 _523_ (.A(net198),
    .TE_B(_097_),
    .Z(la_data_out[36]));
 sky130_fd_sc_hd__ebufn_8 _524_ (.A(net199),
    .TE_B(_098_),
    .Z(la_data_out[37]));
 sky130_fd_sc_hd__ebufn_8 _525_ (.A(net200),
    .TE_B(_099_),
    .Z(la_data_out[38]));
 sky130_fd_sc_hd__ebufn_8 _526_ (.A(net201),
    .TE_B(_100_),
    .Z(la_data_out[39]));
 sky130_fd_sc_hd__ebufn_8 _527_ (.A(net202),
    .TE_B(_101_),
    .Z(la_data_out[40]));
 sky130_fd_sc_hd__ebufn_8 _528_ (.A(net203),
    .TE_B(_102_),
    .Z(la_data_out[41]));
 sky130_fd_sc_hd__ebufn_8 _529_ (.A(net204),
    .TE_B(_103_),
    .Z(la_data_out[42]));
 sky130_fd_sc_hd__ebufn_8 _530_ (.A(net205),
    .TE_B(_104_),
    .Z(la_data_out[43]));
 sky130_fd_sc_hd__ebufn_8 _531_ (.A(net206),
    .TE_B(_105_),
    .Z(la_data_out[44]));
 sky130_fd_sc_hd__ebufn_8 _532_ (.A(net207),
    .TE_B(_106_),
    .Z(la_data_out[45]));
 sky130_fd_sc_hd__ebufn_8 _533_ (.A(net208),
    .TE_B(_107_),
    .Z(la_data_out[46]));
 sky130_fd_sc_hd__ebufn_8 _534_ (.A(net209),
    .TE_B(_108_),
    .Z(la_data_out[47]));
 sky130_fd_sc_hd__ebufn_8 _535_ (.A(net210),
    .TE_B(_109_),
    .Z(la_data_out[48]));
 sky130_fd_sc_hd__ebufn_8 _536_ (.A(net211),
    .TE_B(_110_),
    .Z(la_data_out[49]));
 sky130_fd_sc_hd__ebufn_8 _537_ (.A(net212),
    .TE_B(_111_),
    .Z(la_data_out[50]));
 sky130_fd_sc_hd__ebufn_8 _538_ (.A(net213),
    .TE_B(_112_),
    .Z(la_data_out[51]));
 sky130_fd_sc_hd__ebufn_8 _539_ (.A(net214),
    .TE_B(_113_),
    .Z(la_data_out[52]));
 sky130_fd_sc_hd__ebufn_8 _540_ (.A(net215),
    .TE_B(_114_),
    .Z(la_data_out[53]));
 sky130_fd_sc_hd__ebufn_8 _541_ (.A(net216),
    .TE_B(_115_),
    .Z(la_data_out[54]));
 sky130_fd_sc_hd__ebufn_8 _542_ (.A(net217),
    .TE_B(_116_),
    .Z(la_data_out[55]));
 sky130_fd_sc_hd__ebufn_8 _543_ (.A(net218),
    .TE_B(_117_),
    .Z(la_data_out[56]));
 sky130_fd_sc_hd__ebufn_8 _544_ (.A(net219),
    .TE_B(_118_),
    .Z(la_data_out[57]));
 sky130_fd_sc_hd__ebufn_8 _545_ (.A(net220),
    .TE_B(_119_),
    .Z(la_data_out[58]));
 sky130_fd_sc_hd__ebufn_8 _546_ (.A(net221),
    .TE_B(_120_),
    .Z(la_data_out[59]));
 sky130_fd_sc_hd__ebufn_8 _547_ (.A(net222),
    .TE_B(_121_),
    .Z(la_data_out[60]));
 sky130_fd_sc_hd__ebufn_8 _548_ (.A(net223),
    .TE_B(_122_),
    .Z(la_data_out[61]));
 sky130_fd_sc_hd__ebufn_8 _549_ (.A(net224),
    .TE_B(_123_),
    .Z(la_data_out[62]));
 sky130_fd_sc_hd__ebufn_8 _550_ (.A(net225),
    .TE_B(_124_),
    .Z(la_data_out[63]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_active),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[18]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[19]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(io_in[20]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[21]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[22]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(io_in[23]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(io_in[24]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(io_in[25]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(io_in[26]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(io_in[27]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(io_in[28]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(io_in[29]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(io_in[30]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(io_in[31]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(io_in[32]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(io_in[33]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(io_in[34]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(io_in[35]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(io_in[36]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(io_in[37]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(io_out[9]));
 sky130_fd_sc_hd__conb_1 macro_7_37 (.LO(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__278__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__261__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__259__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__246__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__170__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__159__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_active));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(io_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(io_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(io_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__157__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__286__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__285__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__265__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__284__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__269__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__253__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__236__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__A_N (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__274__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__231__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__A_N (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__B1 (.DIODE(net31));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_624 ();
 assign io_oeb[0] = net226;
 assign io_oeb[10] = net236;
 assign io_oeb[11] = net237;
 assign io_oeb[12] = net238;
 assign io_oeb[13] = net239;
 assign io_oeb[14] = net240;
 assign io_oeb[15] = net241;
 assign io_oeb[16] = net242;
 assign io_oeb[17] = net243;
 assign io_oeb[18] = net244;
 assign io_oeb[19] = net245;
 assign io_oeb[1] = net227;
 assign io_oeb[20] = net246;
 assign io_oeb[21] = net247;
 assign io_oeb[22] = net248;
 assign io_oeb[23] = net249;
 assign io_oeb[24] = net250;
 assign io_oeb[25] = net251;
 assign io_oeb[26] = net252;
 assign io_oeb[27] = net253;
 assign io_oeb[28] = net254;
 assign io_oeb[29] = net255;
 assign io_oeb[2] = net228;
 assign io_oeb[30] = net256;
 assign io_oeb[31] = net257;
 assign io_oeb[32] = net258;
 assign io_oeb[33] = net37;
 assign io_oeb[34] = net38;
 assign io_oeb[35] = net39;
 assign io_oeb[36] = net40;
 assign io_oeb[37] = net41;
 assign io_oeb[3] = net229;
 assign io_oeb[4] = net230;
 assign io_oeb[5] = net231;
 assign io_oeb[6] = net232;
 assign io_oeb[7] = net233;
 assign io_oeb[8] = net234;
 assign io_oeb[9] = net235;
 assign io_out[18] = net45;
 assign io_out[19] = net46;
 assign io_out[1] = net42;
 assign io_out[20] = net47;
 assign io_out[21] = net48;
 assign io_out[22] = net49;
 assign io_out[23] = net50;
 assign io_out[24] = net51;
 assign io_out[25] = net52;
 assign io_out[26] = net53;
 assign io_out[27] = net54;
 assign io_out[28] = net55;
 assign io_out[29] = net56;
 assign io_out[2] = net43;
 assign io_out[30] = net57;
 assign io_out[31] = net58;
 assign io_out[32] = net59;
 assign io_out[33] = net60;
 assign io_out[34] = net61;
 assign io_out[35] = net62;
 assign io_out[36] = net63;
 assign io_out[37] = net64;
 assign io_out[3] = net44;
 assign la_data_out[0] = net65;
 assign la_data_out[100] = net133;
 assign la_data_out[101] = net134;
 assign la_data_out[102] = net135;
 assign la_data_out[103] = net136;
 assign la_data_out[104] = net137;
 assign la_data_out[105] = net138;
 assign la_data_out[106] = net139;
 assign la_data_out[107] = net140;
 assign la_data_out[108] = net141;
 assign la_data_out[109] = net142;
 assign la_data_out[10] = net75;
 assign la_data_out[110] = net143;
 assign la_data_out[111] = net144;
 assign la_data_out[112] = net145;
 assign la_data_out[113] = net146;
 assign la_data_out[114] = net147;
 assign la_data_out[115] = net148;
 assign la_data_out[116] = net149;
 assign la_data_out[117] = net150;
 assign la_data_out[118] = net151;
 assign la_data_out[119] = net152;
 assign la_data_out[11] = net76;
 assign la_data_out[120] = net153;
 assign la_data_out[121] = net154;
 assign la_data_out[122] = net155;
 assign la_data_out[123] = net156;
 assign la_data_out[124] = net157;
 assign la_data_out[125] = net158;
 assign la_data_out[126] = net159;
 assign la_data_out[127] = net160;
 assign la_data_out[12] = net77;
 assign la_data_out[13] = net78;
 assign la_data_out[14] = net79;
 assign la_data_out[15] = net80;
 assign la_data_out[16] = net81;
 assign la_data_out[17] = net82;
 assign la_data_out[18] = net83;
 assign la_data_out[19] = net84;
 assign la_data_out[1] = net66;
 assign la_data_out[20] = net85;
 assign la_data_out[21] = net86;
 assign la_data_out[22] = net87;
 assign la_data_out[23] = net88;
 assign la_data_out[24] = net89;
 assign la_data_out[25] = net90;
 assign la_data_out[26] = net91;
 assign la_data_out[27] = net92;
 assign la_data_out[28] = net93;
 assign la_data_out[29] = net94;
 assign la_data_out[2] = net67;
 assign la_data_out[30] = net95;
 assign la_data_out[31] = net96;
 assign la_data_out[3] = net68;
 assign la_data_out[4] = net69;
 assign la_data_out[5] = net70;
 assign la_data_out[64] = net97;
 assign la_data_out[65] = net98;
 assign la_data_out[66] = net99;
 assign la_data_out[67] = net100;
 assign la_data_out[68] = net101;
 assign la_data_out[69] = net102;
 assign la_data_out[6] = net71;
 assign la_data_out[70] = net103;
 assign la_data_out[71] = net104;
 assign la_data_out[72] = net105;
 assign la_data_out[73] = net106;
 assign la_data_out[74] = net107;
 assign la_data_out[75] = net108;
 assign la_data_out[76] = net109;
 assign la_data_out[77] = net110;
 assign la_data_out[78] = net111;
 assign la_data_out[79] = net112;
 assign la_data_out[7] = net72;
 assign la_data_out[80] = net113;
 assign la_data_out[81] = net114;
 assign la_data_out[82] = net115;
 assign la_data_out[83] = net116;
 assign la_data_out[84] = net117;
 assign la_data_out[85] = net118;
 assign la_data_out[86] = net119;
 assign la_data_out[87] = net120;
 assign la_data_out[88] = net121;
 assign la_data_out[89] = net122;
 assign la_data_out[8] = net73;
 assign la_data_out[90] = net123;
 assign la_data_out[91] = net124;
 assign la_data_out[92] = net125;
 assign la_data_out[93] = net126;
 assign la_data_out[94] = net127;
 assign la_data_out[95] = net128;
 assign la_data_out[96] = net129;
 assign la_data_out[97] = net130;
 assign la_data_out[98] = net131;
 assign la_data_out[99] = net132;
 assign la_data_out[9] = net74;
 assign wbs_ack_o = net161;
 assign wbs_dat_o[0] = net162;
 assign wbs_dat_o[10] = net172;
 assign wbs_dat_o[11] = net173;
 assign wbs_dat_o[12] = net174;
 assign wbs_dat_o[13] = net175;
 assign wbs_dat_o[14] = net176;
 assign wbs_dat_o[15] = net177;
 assign wbs_dat_o[16] = net178;
 assign wbs_dat_o[17] = net179;
 assign wbs_dat_o[18] = net180;
 assign wbs_dat_o[19] = net181;
 assign wbs_dat_o[1] = net163;
 assign wbs_dat_o[20] = net182;
 assign wbs_dat_o[21] = net183;
 assign wbs_dat_o[22] = net184;
 assign wbs_dat_o[23] = net185;
 assign wbs_dat_o[24] = net186;
 assign wbs_dat_o[25] = net187;
 assign wbs_dat_o[26] = net188;
 assign wbs_dat_o[27] = net189;
 assign wbs_dat_o[28] = net190;
 assign wbs_dat_o[29] = net191;
 assign wbs_dat_o[2] = net164;
 assign wbs_dat_o[30] = net192;
 assign wbs_dat_o[31] = net193;
 assign wbs_dat_o[3] = net165;
 assign wbs_dat_o[4] = net166;
 assign wbs_dat_o[5] = net167;
 assign wbs_dat_o[6] = net168;
 assign wbs_dat_o[7] = net169;
 assign wbs_dat_o[8] = net170;
 assign wbs_dat_o[9] = net171;
endmodule

