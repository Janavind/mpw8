// This is the unpowered netlist.
module macro_decap_3 (io_active,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input io_active;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net228;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net229;
 wire net257;
 wire net258;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net46;
 wire net47;
 wire net43;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net44;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net45;
 wire net66;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net76;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net77;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net67;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net68;
 wire net96;
 wire net97;
 wire net69;
 wire net70;
 wire net71;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net72;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net73;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net74;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net75;
 wire net162;
 wire net163;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net164;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net165;
 wire net193;
 wire net194;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;

 sky130_fd_sc_hd__inv_2 _157_ (.A(net1),
    .Y(_124_));
 sky130_fd_sc_hd__buf_4 _158_ (.A(net1),
    .X(_089_));
 sky130_fd_sc_hd__buf_4 _159_ (.A(_089_),
    .X(_090_));
 sky130_fd_sc_hd__inv_2 _160_ (.A(_090_),
    .Y(_123_));
 sky130_fd_sc_hd__inv_2 _161_ (.A(_090_),
    .Y(_122_));
 sky130_fd_sc_hd__inv_2 _162_ (.A(_090_),
    .Y(_121_));
 sky130_fd_sc_hd__inv_2 _163_ (.A(_090_),
    .Y(_120_));
 sky130_fd_sc_hd__inv_2 _164_ (.A(_090_),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _165_ (.A(_090_),
    .Y(_118_));
 sky130_fd_sc_hd__inv_2 _166_ (.A(_090_),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _167_ (.A(_090_),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _168_ (.A(_090_),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _169_ (.A(_090_),
    .Y(_114_));
 sky130_fd_sc_hd__buf_4 _170_ (.A(_089_),
    .X(_091_));
 sky130_fd_sc_hd__inv_2 _171_ (.A(_091_),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _172_ (.A(_091_),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _173_ (.A(_091_),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _174_ (.A(_091_),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _175_ (.A(_091_),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _176_ (.A(_091_),
    .Y(_108_));
 sky130_fd_sc_hd__inv_2 _177_ (.A(_091_),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _178_ (.A(_091_),
    .Y(_106_));
 sky130_fd_sc_hd__inv_2 _179_ (.A(_091_),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _180_ (.A(_091_),
    .Y(_104_));
 sky130_fd_sc_hd__buf_4 _181_ (.A(_089_),
    .X(_092_));
 sky130_fd_sc_hd__inv_2 _182_ (.A(_092_),
    .Y(_103_));
 sky130_fd_sc_hd__inv_2 _183_ (.A(_092_),
    .Y(_102_));
 sky130_fd_sc_hd__inv_2 _184_ (.A(_092_),
    .Y(_101_));
 sky130_fd_sc_hd__inv_2 _185_ (.A(_092_),
    .Y(_100_));
 sky130_fd_sc_hd__inv_2 _186_ (.A(_092_),
    .Y(_099_));
 sky130_fd_sc_hd__inv_2 _187_ (.A(_092_),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _188_ (.A(_092_),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _189_ (.A(_092_),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _190_ (.A(_092_),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _191_ (.A(_092_),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _192_ (.A(_089_),
    .Y(_093_));
 sky130_fd_sc_hd__nand2b_1 _193_ (.A_N(net19),
    .B(net18),
    .Y(_000_));
 sky130_fd_sc_hd__o31a_1 _194_ (.A1(net8),
    .A2(net6),
    .A3(net7),
    .B1(_000_),
    .X(_001_));
 sky130_fd_sc_hd__xnor2_1 _195_ (.A(net9),
    .B(_001_),
    .Y(_002_));
 sky130_fd_sc_hd__or2_1 _196_ (.A(net5),
    .B(_002_),
    .X(_003_));
 sky130_fd_sc_hd__o21a_1 _197_ (.A1(net6),
    .A2(net7),
    .B1(_000_),
    .X(_004_));
 sky130_fd_sc_hd__xnor2_1 _198_ (.A(net8),
    .B(_004_),
    .Y(_005_));
 sky130_fd_sc_hd__or2_1 _199_ (.A(net4),
    .B(_005_),
    .X(_006_));
 sky130_fd_sc_hd__nand3b_1 _200_ (.A_N(net7),
    .B(_000_),
    .C(net6),
    .Y(_007_));
 sky130_fd_sc_hd__a21bo_1 _201_ (.A1(net6),
    .A2(_000_),
    .B1_N(net7),
    .X(_008_));
 sky130_fd_sc_hd__a21o_1 _202_ (.A1(_007_),
    .A2(_008_),
    .B1(net3),
    .X(_009_));
 sky130_fd_sc_hd__or2b_1 _203_ (.A(net2),
    .B_N(net6),
    .X(_010_));
 sky130_fd_sc_hd__and3_1 _204_ (.A(net3),
    .B(_007_),
    .C(_008_),
    .X(_011_));
 sky130_fd_sc_hd__a21o_1 _205_ (.A1(_009_),
    .A2(_010_),
    .B1(_011_),
    .X(_012_));
 sky130_fd_sc_hd__and2_1 _206_ (.A(net5),
    .B(_002_),
    .X(_013_));
 sky130_fd_sc_hd__and2_1 _207_ (.A(net4),
    .B(_005_),
    .X(_014_));
 sky130_fd_sc_hd__a211o_1 _208_ (.A1(_006_),
    .A2(_012_),
    .B1(_013_),
    .C1(_014_),
    .X(_015_));
 sky130_fd_sc_hd__a21oi_1 _209_ (.A1(net9),
    .A2(_000_),
    .B1(_001_),
    .Y(_016_));
 sky130_fd_sc_hd__a21oi_1 _210_ (.A1(_003_),
    .A2(_015_),
    .B1(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__a31o_1 _211_ (.A1(_016_),
    .A2(_003_),
    .A3(_015_),
    .B1(net19),
    .X(_018_));
 sky130_fd_sc_hd__or2_1 _212_ (.A(_017_),
    .B(_018_),
    .X(_019_));
 sky130_fd_sc_hd__nand2b_1 _213_ (.A_N(net21),
    .B(net20),
    .Y(_020_));
 sky130_fd_sc_hd__o31a_1 _214_ (.A1(net16),
    .A2(net14),
    .A3(net15),
    .B1(_020_),
    .X(_021_));
 sky130_fd_sc_hd__xnor2_1 _215_ (.A(net17),
    .B(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__or2_1 _216_ (.A(net13),
    .B(_022_),
    .X(_023_));
 sky130_fd_sc_hd__o21a_1 _217_ (.A1(net14),
    .A2(net15),
    .B1(_020_),
    .X(_024_));
 sky130_fd_sc_hd__xnor2_1 _218_ (.A(net16),
    .B(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__or2_1 _219_ (.A(net12),
    .B(_025_),
    .X(_026_));
 sky130_fd_sc_hd__nand3b_1 _220_ (.A_N(net15),
    .B(_020_),
    .C(net14),
    .Y(_027_));
 sky130_fd_sc_hd__a21bo_1 _221_ (.A1(net14),
    .A2(_020_),
    .B1_N(net15),
    .X(_028_));
 sky130_fd_sc_hd__a21o_1 _222_ (.A1(_027_),
    .A2(_028_),
    .B1(net11),
    .X(_029_));
 sky130_fd_sc_hd__or2b_1 _223_ (.A(net10),
    .B_N(net14),
    .X(_030_));
 sky130_fd_sc_hd__and3_1 _224_ (.A(net11),
    .B(_027_),
    .C(_028_),
    .X(_031_));
 sky130_fd_sc_hd__a21o_1 _225_ (.A1(_029_),
    .A2(_030_),
    .B1(_031_),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _226_ (.A(net13),
    .B(_022_),
    .X(_033_));
 sky130_fd_sc_hd__and2_1 _227_ (.A(net12),
    .B(_025_),
    .X(_034_));
 sky130_fd_sc_hd__a211o_1 _228_ (.A1(_026_),
    .A2(_032_),
    .B1(_033_),
    .C1(_034_),
    .X(_035_));
 sky130_fd_sc_hd__a21oi_1 _229_ (.A1(net17),
    .A2(_020_),
    .B1(_021_),
    .Y(_036_));
 sky130_fd_sc_hd__a21oi_1 _230_ (.A1(_023_),
    .A2(_035_),
    .B1(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__a31o_1 _231_ (.A1(_036_),
    .A2(_023_),
    .A3(_035_),
    .B1(net21),
    .X(_038_));
 sky130_fd_sc_hd__or2_1 _232_ (.A(_037_),
    .B(_038_),
    .X(_039_));
 sky130_fd_sc_hd__nor3_2 _233_ (.A(_124_),
    .B(_037_),
    .C(_038_),
    .Y(net31));
 sky130_fd_sc_hd__nor3_1 _234_ (.A(_124_),
    .B(_017_),
    .C(_018_),
    .Y(net32));
 sky130_fd_sc_hd__o22a_1 _235_ (.A1(_019_),
    .A2(_039_),
    .B1(net31),
    .B2(net32),
    .X(net22));
 sky130_fd_sc_hd__inv_2 _236_ (.A(net19),
    .Y(_040_));
 sky130_fd_sc_hd__o2bb2a_1 _237_ (.A1_N(net6),
    .A2_N(net2),
    .B1(_040_),
    .B2(net18),
    .X(_041_));
 sky130_fd_sc_hd__o21a_1 _238_ (.A1(net6),
    .A2(net2),
    .B1(_041_),
    .X(_042_));
 sky130_fd_sc_hd__a31o_1 _239_ (.A1(net6),
    .A2(net19),
    .A3(net2),
    .B1(_042_),
    .X(_043_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(net21),
    .Y(_044_));
 sky130_fd_sc_hd__o2bb2a_1 _241_ (.A1_N(net14),
    .A2_N(net10),
    .B1(_044_),
    .B2(net20),
    .X(_045_));
 sky130_fd_sc_hd__o21a_1 _242_ (.A1(net14),
    .A2(net10),
    .B1(_045_),
    .X(_046_));
 sky130_fd_sc_hd__a31o_1 _243_ (.A1(net14),
    .A2(net21),
    .A3(net10),
    .B1(_046_),
    .X(_047_));
 sky130_fd_sc_hd__and2_1 _244_ (.A(_089_),
    .B(_047_),
    .X(_048_));
 sky130_fd_sc_hd__clkbuf_1 _245_ (.A(_048_),
    .X(net23));
 sky130_fd_sc_hd__and2_1 _246_ (.A(_089_),
    .B(_043_),
    .X(_049_));
 sky130_fd_sc_hd__clkbuf_1 _247_ (.A(_049_),
    .X(net27));
 sky130_fd_sc_hd__o2bb2a_1 _248_ (.A1_N(_043_),
    .A2_N(_047_),
    .B1(net23),
    .B2(net27),
    .X(net33));
 sky130_fd_sc_hd__or2b_1 _249_ (.A(_011_),
    .B_N(_009_),
    .X(_050_));
 sky130_fd_sc_hd__xnor2_1 _250_ (.A(_050_),
    .B(_010_),
    .Y(_051_));
 sky130_fd_sc_hd__o21a_1 _251_ (.A1(net7),
    .A2(net18),
    .B1(net3),
    .X(_052_));
 sky130_fd_sc_hd__a211o_1 _252_ (.A1(net7),
    .A2(net18),
    .B1(_040_),
    .C1(_052_),
    .X(_053_));
 sky130_fd_sc_hd__o21a_1 _253_ (.A1(net19),
    .A2(_051_),
    .B1(_053_),
    .X(_054_));
 sky130_fd_sc_hd__or2b_1 _254_ (.A(_031_),
    .B_N(_029_),
    .X(_055_));
 sky130_fd_sc_hd__xnor2_1 _255_ (.A(_055_),
    .B(_030_),
    .Y(_056_));
 sky130_fd_sc_hd__o21a_1 _256_ (.A1(net15),
    .A2(net20),
    .B1(net11),
    .X(_057_));
 sky130_fd_sc_hd__a211o_1 _257_ (.A1(net15),
    .A2(net20),
    .B1(_044_),
    .C1(_057_),
    .X(_058_));
 sky130_fd_sc_hd__o21a_1 _258_ (.A1(net21),
    .A2(_056_),
    .B1(_058_),
    .X(_059_));
 sky130_fd_sc_hd__and2_1 _259_ (.A(_089_),
    .B(_059_),
    .X(_060_));
 sky130_fd_sc_hd__clkbuf_1 _260_ (.A(_060_),
    .X(net24));
 sky130_fd_sc_hd__and2_1 _261_ (.A(_089_),
    .B(_054_),
    .X(_061_));
 sky130_fd_sc_hd__clkbuf_1 _262_ (.A(_061_),
    .X(net28));
 sky130_fd_sc_hd__o2bb2a_1 _263_ (.A1_N(_054_),
    .A2_N(_059_),
    .B1(net24),
    .B2(net28),
    .X(net34));
 sky130_fd_sc_hd__a21o_1 _264_ (.A1(net18),
    .A2(net4),
    .B1(net8),
    .X(_062_));
 sky130_fd_sc_hd__or2_1 _265_ (.A(net18),
    .B(net4),
    .X(_063_));
 sky130_fd_sc_hd__xor2_1 _266_ (.A(net4),
    .B(_005_),
    .X(_064_));
 sky130_fd_sc_hd__or2_1 _267_ (.A(_064_),
    .B(_012_),
    .X(_065_));
 sky130_fd_sc_hd__a21oi_1 _268_ (.A1(_064_),
    .A2(_012_),
    .B1(net19),
    .Y(_066_));
 sky130_fd_sc_hd__a32o_1 _269_ (.A1(net19),
    .A2(_062_),
    .A3(_063_),
    .B1(_065_),
    .B2(_066_),
    .X(_067_));
 sky130_fd_sc_hd__a21o_1 _270_ (.A1(net20),
    .A2(net12),
    .B1(net16),
    .X(_068_));
 sky130_fd_sc_hd__or2_1 _271_ (.A(net20),
    .B(net12),
    .X(_069_));
 sky130_fd_sc_hd__xor2_1 _272_ (.A(net12),
    .B(_025_),
    .X(_070_));
 sky130_fd_sc_hd__or2_1 _273_ (.A(_070_),
    .B(_032_),
    .X(_071_));
 sky130_fd_sc_hd__a21oi_1 _274_ (.A1(_070_),
    .A2(_032_),
    .B1(net21),
    .Y(_072_));
 sky130_fd_sc_hd__a32o_1 _275_ (.A1(net21),
    .A2(_068_),
    .A3(_069_),
    .B1(_071_),
    .B2(_072_),
    .X(_073_));
 sky130_fd_sc_hd__and2_1 _276_ (.A(net1),
    .B(_073_),
    .X(_074_));
 sky130_fd_sc_hd__clkbuf_1 _277_ (.A(_074_),
    .X(net25));
 sky130_fd_sc_hd__and2_1 _278_ (.A(_089_),
    .B(_067_),
    .X(_075_));
 sky130_fd_sc_hd__clkbuf_1 _279_ (.A(_075_),
    .X(net29));
 sky130_fd_sc_hd__o2bb2a_1 _280_ (.A1_N(_067_),
    .A2_N(_073_),
    .B1(net25),
    .B2(net29),
    .X(net35));
 sky130_fd_sc_hd__a21oi_1 _281_ (.A1(_006_),
    .A2(_012_),
    .B1(_014_),
    .Y(_076_));
 sky130_fd_sc_hd__and2b_1 _282_ (.A_N(_013_),
    .B(_003_),
    .X(_077_));
 sky130_fd_sc_hd__xnor2_1 _283_ (.A(_076_),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__nor2_1 _284_ (.A(net19),
    .B(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__o21a_1 _285_ (.A1(net9),
    .A2(net18),
    .B1(net5),
    .X(_080_));
 sky130_fd_sc_hd__a21o_1 _286_ (.A1(net9),
    .A2(net18),
    .B1(_040_),
    .X(_081_));
 sky130_fd_sc_hd__nor2_1 _287_ (.A(_080_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__a21o_1 _288_ (.A1(_026_),
    .A2(_032_),
    .B1(_034_),
    .X(_083_));
 sky130_fd_sc_hd__and2b_1 _289_ (.A_N(_033_),
    .B(_023_),
    .X(_084_));
 sky130_fd_sc_hd__xnor2_1 _290_ (.A(_083_),
    .B(_084_),
    .Y(_085_));
 sky130_fd_sc_hd__o21a_1 _291_ (.A1(net17),
    .A2(net20),
    .B1(net13),
    .X(_086_));
 sky130_fd_sc_hd__a211oi_2 _292_ (.A1(net17),
    .A2(net20),
    .B1(_044_),
    .C1(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__a21o_1 _293_ (.A1(_044_),
    .A2(_085_),
    .B1(_087_),
    .X(_088_));
 sky130_fd_sc_hd__a211oi_2 _294_ (.A1(_044_),
    .A2(_085_),
    .B1(_087_),
    .C1(_124_),
    .Y(net26));
 sky130_fd_sc_hd__o221a_1 _295_ (.A1(net19),
    .A2(_078_),
    .B1(_080_),
    .B2(_081_),
    .C1(_089_),
    .X(net30));
 sky130_fd_sc_hd__o32a_1 _296_ (.A1(_079_),
    .A2(_082_),
    .A3(_088_),
    .B1(net26),
    .B2(net30),
    .X(net36));
 sky130_fd_sc_hd__conb_1 macro_decap_3_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 macro_decap_3_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 macro_decap_3_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 macro_decap_3_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 macro_decap_3_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 macro_decap_3_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 macro_decap_3_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 macro_decap_3_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 macro_decap_3_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 macro_decap_3_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 macro_decap_3_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 macro_decap_3_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 macro_decap_3_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 macro_decap_3_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 macro_decap_3_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 macro_decap_3_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 macro_decap_3_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 macro_decap_3_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 macro_decap_3_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 macro_decap_3_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 macro_decap_3_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 macro_decap_3_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 macro_decap_3_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 macro_decap_3_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 macro_decap_3_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 macro_decap_3_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 macro_decap_3_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 macro_decap_3_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 macro_decap_3_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 macro_decap_3_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 macro_decap_3_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 macro_decap_3_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 macro_decap_3_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 macro_decap_3_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 macro_decap_3_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 macro_decap_3_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 macro_decap_3_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 macro_decap_3_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 macro_decap_3_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 macro_decap_3_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 macro_decap_3_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 macro_decap_3_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 macro_decap_3_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 macro_decap_3_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 macro_decap_3_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 macro_decap_3_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 macro_decap_3_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 macro_decap_3_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 macro_decap_3_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 macro_decap_3_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 macro_decap_3_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 macro_decap_3_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 macro_decap_3_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 macro_decap_3_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 macro_decap_3_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 macro_decap_3_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 macro_decap_3_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 macro_decap_3_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 macro_decap_3_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 macro_decap_3_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 macro_decap_3_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 macro_decap_3_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 macro_decap_3_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 macro_decap_3_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 macro_decap_3_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 macro_decap_3_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 macro_decap_3_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 macro_decap_3_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 macro_decap_3_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 macro_decap_3_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 macro_decap_3_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 macro_decap_3_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 macro_decap_3_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 macro_decap_3_111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 macro_decap_3_112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 macro_decap_3_113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 macro_decap_3_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 macro_decap_3_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 macro_decap_3_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 macro_decap_3_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 macro_decap_3_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 macro_decap_3_119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 macro_decap_3_120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 macro_decap_3_121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 macro_decap_3_122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 macro_decap_3_123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 macro_decap_3_124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 macro_decap_3_125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 macro_decap_3_126 (.LO(net126));
 sky130_fd_sc_hd__conb_1 macro_decap_3_127 (.LO(net127));
 sky130_fd_sc_hd__conb_1 macro_decap_3_128 (.LO(net128));
 sky130_fd_sc_hd__conb_1 macro_decap_3_129 (.LO(net129));
 sky130_fd_sc_hd__conb_1 macro_decap_3_130 (.LO(net130));
 sky130_fd_sc_hd__conb_1 macro_decap_3_131 (.LO(net131));
 sky130_fd_sc_hd__conb_1 macro_decap_3_132 (.LO(net132));
 sky130_fd_sc_hd__conb_1 macro_decap_3_133 (.LO(net133));
 sky130_fd_sc_hd__conb_1 macro_decap_3_134 (.LO(net134));
 sky130_fd_sc_hd__conb_1 macro_decap_3_135 (.LO(net135));
 sky130_fd_sc_hd__conb_1 macro_decap_3_136 (.LO(net136));
 sky130_fd_sc_hd__conb_1 macro_decap_3_137 (.LO(net137));
 sky130_fd_sc_hd__conb_1 macro_decap_3_138 (.LO(net138));
 sky130_fd_sc_hd__conb_1 macro_decap_3_139 (.LO(net139));
 sky130_fd_sc_hd__conb_1 macro_decap_3_140 (.LO(net140));
 sky130_fd_sc_hd__conb_1 macro_decap_3_141 (.LO(net141));
 sky130_fd_sc_hd__conb_1 macro_decap_3_142 (.LO(net142));
 sky130_fd_sc_hd__conb_1 macro_decap_3_143 (.LO(net143));
 sky130_fd_sc_hd__conb_1 macro_decap_3_144 (.LO(net144));
 sky130_fd_sc_hd__conb_1 macro_decap_3_145 (.LO(net145));
 sky130_fd_sc_hd__conb_1 macro_decap_3_146 (.LO(net146));
 sky130_fd_sc_hd__conb_1 macro_decap_3_147 (.LO(net147));
 sky130_fd_sc_hd__conb_1 macro_decap_3_148 (.LO(net148));
 sky130_fd_sc_hd__conb_1 macro_decap_3_149 (.LO(net149));
 sky130_fd_sc_hd__conb_1 macro_decap_3_150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 macro_decap_3_151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 macro_decap_3_152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 macro_decap_3_153 (.LO(net153));
 sky130_fd_sc_hd__conb_1 macro_decap_3_154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 macro_decap_3_155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 macro_decap_3_156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 macro_decap_3_157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 macro_decap_3_158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 macro_decap_3_159 (.LO(net159));
 sky130_fd_sc_hd__conb_1 macro_decap_3_160 (.LO(net160));
 sky130_fd_sc_hd__conb_1 macro_decap_3_161 (.LO(net161));
 sky130_fd_sc_hd__conb_1 macro_decap_3_162 (.LO(net162));
 sky130_fd_sc_hd__conb_1 macro_decap_3_163 (.LO(net163));
 sky130_fd_sc_hd__conb_1 macro_decap_3_164 (.LO(net164));
 sky130_fd_sc_hd__conb_1 macro_decap_3_165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 macro_decap_3_166 (.LO(net166));
 sky130_fd_sc_hd__conb_1 macro_decap_3_167 (.LO(net167));
 sky130_fd_sc_hd__conb_1 macro_decap_3_168 (.LO(net168));
 sky130_fd_sc_hd__conb_1 macro_decap_3_169 (.LO(net169));
 sky130_fd_sc_hd__conb_1 macro_decap_3_170 (.LO(net170));
 sky130_fd_sc_hd__conb_1 macro_decap_3_171 (.LO(net171));
 sky130_fd_sc_hd__conb_1 macro_decap_3_172 (.LO(net172));
 sky130_fd_sc_hd__conb_1 macro_decap_3_173 (.LO(net173));
 sky130_fd_sc_hd__conb_1 macro_decap_3_174 (.LO(net174));
 sky130_fd_sc_hd__conb_1 macro_decap_3_175 (.LO(net175));
 sky130_fd_sc_hd__conb_1 macro_decap_3_176 (.LO(net176));
 sky130_fd_sc_hd__conb_1 macro_decap_3_177 (.LO(net177));
 sky130_fd_sc_hd__conb_1 macro_decap_3_178 (.LO(net178));
 sky130_fd_sc_hd__conb_1 macro_decap_3_179 (.LO(net179));
 sky130_fd_sc_hd__conb_1 macro_decap_3_180 (.LO(net180));
 sky130_fd_sc_hd__conb_1 macro_decap_3_181 (.LO(net181));
 sky130_fd_sc_hd__conb_1 macro_decap_3_182 (.LO(net182));
 sky130_fd_sc_hd__conb_1 macro_decap_3_183 (.LO(net183));
 sky130_fd_sc_hd__conb_1 macro_decap_3_184 (.LO(net184));
 sky130_fd_sc_hd__conb_1 macro_decap_3_185 (.LO(net185));
 sky130_fd_sc_hd__conb_1 macro_decap_3_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 macro_decap_3_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 macro_decap_3_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 macro_decap_3_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 macro_decap_3_190 (.LO(net190));
 sky130_fd_sc_hd__conb_1 macro_decap_3_191 (.LO(net191));
 sky130_fd_sc_hd__conb_1 macro_decap_3_192 (.LO(net192));
 sky130_fd_sc_hd__conb_1 macro_decap_3_193 (.LO(net193));
 sky130_fd_sc_hd__conb_1 _519__194 (.LO(net194));
 sky130_fd_sc_hd__conb_1 _520__195 (.LO(net195));
 sky130_fd_sc_hd__conb_1 _521__196 (.LO(net196));
 sky130_fd_sc_hd__conb_1 _522__197 (.LO(net197));
 sky130_fd_sc_hd__conb_1 _523__198 (.LO(net198));
 sky130_fd_sc_hd__conb_1 _524__199 (.LO(net199));
 sky130_fd_sc_hd__conb_1 _525__200 (.LO(net200));
 sky130_fd_sc_hd__conb_1 _526__201 (.LO(net201));
 sky130_fd_sc_hd__conb_1 _527__202 (.LO(net202));
 sky130_fd_sc_hd__conb_1 _528__203 (.LO(net203));
 sky130_fd_sc_hd__conb_1 _529__204 (.LO(net204));
 sky130_fd_sc_hd__conb_1 _530__205 (.LO(net205));
 sky130_fd_sc_hd__conb_1 _531__206 (.LO(net206));
 sky130_fd_sc_hd__conb_1 _532__207 (.LO(net207));
 sky130_fd_sc_hd__conb_1 _533__208 (.LO(net208));
 sky130_fd_sc_hd__conb_1 _534__209 (.LO(net209));
 sky130_fd_sc_hd__conb_1 _535__210 (.LO(net210));
 sky130_fd_sc_hd__conb_1 _536__211 (.LO(net211));
 sky130_fd_sc_hd__conb_1 _537__212 (.LO(net212));
 sky130_fd_sc_hd__conb_1 _538__213 (.LO(net213));
 sky130_fd_sc_hd__conb_1 _539__214 (.LO(net214));
 sky130_fd_sc_hd__conb_1 _540__215 (.LO(net215));
 sky130_fd_sc_hd__conb_1 _541__216 (.LO(net216));
 sky130_fd_sc_hd__conb_1 _542__217 (.LO(net217));
 sky130_fd_sc_hd__conb_1 _543__218 (.LO(net218));
 sky130_fd_sc_hd__conb_1 _544__219 (.LO(net219));
 sky130_fd_sc_hd__conb_1 _545__220 (.LO(net220));
 sky130_fd_sc_hd__conb_1 _546__221 (.LO(net221));
 sky130_fd_sc_hd__conb_1 _547__222 (.LO(net222));
 sky130_fd_sc_hd__conb_1 _548__223 (.LO(net223));
 sky130_fd_sc_hd__conb_1 _549__224 (.LO(net224));
 sky130_fd_sc_hd__conb_1 _550__225 (.LO(net225));
 sky130_fd_sc_hd__conb_1 macro_decap_3_226 (.LO(net226));
 sky130_fd_sc_hd__conb_1 macro_decap_3_227 (.LO(net227));
 sky130_fd_sc_hd__conb_1 macro_decap_3_228 (.LO(net228));
 sky130_fd_sc_hd__conb_1 macro_decap_3_229 (.LO(net229));
 sky130_fd_sc_hd__conb_1 macro_decap_3_230 (.LO(net230));
 sky130_fd_sc_hd__conb_1 macro_decap_3_231 (.LO(net231));
 sky130_fd_sc_hd__conb_1 macro_decap_3_232 (.LO(net232));
 sky130_fd_sc_hd__conb_1 macro_decap_3_233 (.LO(net233));
 sky130_fd_sc_hd__conb_1 macro_decap_3_234 (.LO(net234));
 sky130_fd_sc_hd__conb_1 macro_decap_3_235 (.LO(net235));
 sky130_fd_sc_hd__conb_1 macro_decap_3_236 (.LO(net236));
 sky130_fd_sc_hd__conb_1 macro_decap_3_237 (.LO(net237));
 sky130_fd_sc_hd__conb_1 macro_decap_3_238 (.LO(net238));
 sky130_fd_sc_hd__conb_1 macro_decap_3_239 (.LO(net239));
 sky130_fd_sc_hd__conb_1 macro_decap_3_240 (.LO(net240));
 sky130_fd_sc_hd__conb_1 macro_decap_3_241 (.LO(net241));
 sky130_fd_sc_hd__conb_1 macro_decap_3_242 (.LO(net242));
 sky130_fd_sc_hd__conb_1 macro_decap_3_243 (.LO(net243));
 sky130_fd_sc_hd__conb_1 macro_decap_3_244 (.LO(net244));
 sky130_fd_sc_hd__conb_1 macro_decap_3_245 (.LO(net245));
 sky130_fd_sc_hd__conb_1 macro_decap_3_246 (.LO(net246));
 sky130_fd_sc_hd__conb_1 macro_decap_3_247 (.LO(net247));
 sky130_fd_sc_hd__conb_1 macro_decap_3_248 (.LO(net248));
 sky130_fd_sc_hd__conb_1 macro_decap_3_249 (.LO(net249));
 sky130_fd_sc_hd__conb_1 macro_decap_3_250 (.LO(net250));
 sky130_fd_sc_hd__conb_1 macro_decap_3_251 (.LO(net251));
 sky130_fd_sc_hd__conb_1 macro_decap_3_252 (.LO(net252));
 sky130_fd_sc_hd__conb_1 macro_decap_3_253 (.LO(net253));
 sky130_fd_sc_hd__conb_1 macro_decap_3_254 (.LO(net254));
 sky130_fd_sc_hd__conb_1 macro_decap_3_255 (.LO(net255));
 sky130_fd_sc_hd__conb_1 macro_decap_3_256 (.LO(net256));
 sky130_fd_sc_hd__conb_1 macro_decap_3_257 (.LO(net257));
 sky130_fd_sc_hd__conb_1 macro_decap_3_258 (.LO(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__C1 (.DIODE(_089_));
 sky130_fd_sc_hd__ebufn_8 _519_ (.A(net194),
    .TE_B(_093_),
    .Z(la_data_out[32]));
 sky130_fd_sc_hd__ebufn_8 _520_ (.A(net195),
    .TE_B(_094_),
    .Z(la_data_out[33]));
 sky130_fd_sc_hd__ebufn_8 _521_ (.A(net196),
    .TE_B(_095_),
    .Z(la_data_out[34]));
 sky130_fd_sc_hd__ebufn_8 _522_ (.A(net197),
    .TE_B(_096_),
    .Z(la_data_out[35]));
 sky130_fd_sc_hd__ebufn_8 _523_ (.A(net198),
    .TE_B(_097_),
    .Z(la_data_out[36]));
 sky130_fd_sc_hd__ebufn_8 _524_ (.A(net199),
    .TE_B(_098_),
    .Z(la_data_out[37]));
 sky130_fd_sc_hd__ebufn_8 _525_ (.A(net200),
    .TE_B(_099_),
    .Z(la_data_out[38]));
 sky130_fd_sc_hd__ebufn_8 _526_ (.A(net201),
    .TE_B(_100_),
    .Z(la_data_out[39]));
 sky130_fd_sc_hd__ebufn_8 _527_ (.A(net202),
    .TE_B(_101_),
    .Z(la_data_out[40]));
 sky130_fd_sc_hd__ebufn_8 _528_ (.A(net203),
    .TE_B(_102_),
    .Z(la_data_out[41]));
 sky130_fd_sc_hd__ebufn_8 _529_ (.A(net204),
    .TE_B(_103_),
    .Z(la_data_out[42]));
 sky130_fd_sc_hd__ebufn_8 _530_ (.A(net205),
    .TE_B(_104_),
    .Z(la_data_out[43]));
 sky130_fd_sc_hd__ebufn_8 _531_ (.A(net206),
    .TE_B(_105_),
    .Z(la_data_out[44]));
 sky130_fd_sc_hd__ebufn_8 _532_ (.A(net207),
    .TE_B(_106_),
    .Z(la_data_out[45]));
 sky130_fd_sc_hd__ebufn_8 _533_ (.A(net208),
    .TE_B(_107_),
    .Z(la_data_out[46]));
 sky130_fd_sc_hd__ebufn_8 _534_ (.A(net209),
    .TE_B(_108_),
    .Z(la_data_out[47]));
 sky130_fd_sc_hd__ebufn_8 _535_ (.A(net210),
    .TE_B(_109_),
    .Z(la_data_out[48]));
 sky130_fd_sc_hd__ebufn_8 _536_ (.A(net211),
    .TE_B(_110_),
    .Z(la_data_out[49]));
 sky130_fd_sc_hd__ebufn_8 _537_ (.A(net212),
    .TE_B(_111_),
    .Z(la_data_out[50]));
 sky130_fd_sc_hd__ebufn_8 _538_ (.A(net213),
    .TE_B(_112_),
    .Z(la_data_out[51]));
 sky130_fd_sc_hd__ebufn_8 _539_ (.A(net214),
    .TE_B(_113_),
    .Z(la_data_out[52]));
 sky130_fd_sc_hd__ebufn_8 _540_ (.A(net215),
    .TE_B(_114_),
    .Z(la_data_out[53]));
 sky130_fd_sc_hd__ebufn_8 _541_ (.A(net216),
    .TE_B(_115_),
    .Z(la_data_out[54]));
 sky130_fd_sc_hd__ebufn_8 _542_ (.A(net217),
    .TE_B(_116_),
    .Z(la_data_out[55]));
 sky130_fd_sc_hd__ebufn_8 _543_ (.A(net218),
    .TE_B(_117_),
    .Z(la_data_out[56]));
 sky130_fd_sc_hd__ebufn_8 _544_ (.A(net219),
    .TE_B(_118_),
    .Z(la_data_out[57]));
 sky130_fd_sc_hd__ebufn_8 _545_ (.A(net220),
    .TE_B(_119_),
    .Z(la_data_out[58]));
 sky130_fd_sc_hd__ebufn_8 _546_ (.A(net221),
    .TE_B(_120_),
    .Z(la_data_out[59]));
 sky130_fd_sc_hd__ebufn_8 _547_ (.A(net222),
    .TE_B(_121_),
    .Z(la_data_out[60]));
 sky130_fd_sc_hd__ebufn_8 _548_ (.A(net223),
    .TE_B(_122_),
    .Z(la_data_out[61]));
 sky130_fd_sc_hd__ebufn_8 _549_ (.A(net224),
    .TE_B(_123_),
    .Z(la_data_out[62]));
 sky130_fd_sc_hd__ebufn_8 _550_ (.A(net225),
    .TE_B(_124_),
    .Z(la_data_out[63]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_active),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[18]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[19]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(io_in[20]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[21]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[22]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(io_in[23]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(io_in[24]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(io_in[25]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(io_in[26]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(io_in[27]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(io_in[28]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(io_in[29]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(io_in[30]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(io_in[31]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(io_in[32]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(io_in[33]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(io_in[34]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(io_in[35]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(io_in[36]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(io_in[37]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(io_out[9]));
 sky130_fd_sc_hd__conb_1 macro_decap_3_37 (.LO(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__278__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__261__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__259__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__246__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__170__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__159__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_active));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(io_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(io_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(io_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__157__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__286__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__285__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__265__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__284__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__269__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__253__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__236__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__A_N (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__274__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__231__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__A_N (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__B1 (.DIODE(net31));
 sky130_fd_sc_hd__fill_8 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_150 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_492 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_456 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_413 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_400 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_57 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_617 ();
 assign io_oeb[0] = net226;
 assign io_oeb[10] = net236;
 assign io_oeb[11] = net237;
 assign io_oeb[12] = net238;
 assign io_oeb[13] = net239;
 assign io_oeb[14] = net240;
 assign io_oeb[15] = net241;
 assign io_oeb[16] = net242;
 assign io_oeb[17] = net243;
 assign io_oeb[18] = net244;
 assign io_oeb[19] = net245;
 assign io_oeb[1] = net227;
 assign io_oeb[20] = net246;
 assign io_oeb[21] = net247;
 assign io_oeb[22] = net248;
 assign io_oeb[23] = net249;
 assign io_oeb[24] = net250;
 assign io_oeb[25] = net251;
 assign io_oeb[26] = net252;
 assign io_oeb[27] = net253;
 assign io_oeb[28] = net254;
 assign io_oeb[29] = net255;
 assign io_oeb[2] = net228;
 assign io_oeb[30] = net256;
 assign io_oeb[31] = net257;
 assign io_oeb[32] = net258;
 assign io_oeb[33] = net37;
 assign io_oeb[34] = net38;
 assign io_oeb[35] = net39;
 assign io_oeb[36] = net40;
 assign io_oeb[37] = net41;
 assign io_oeb[3] = net229;
 assign io_oeb[4] = net230;
 assign io_oeb[5] = net231;
 assign io_oeb[6] = net232;
 assign io_oeb[7] = net233;
 assign io_oeb[8] = net234;
 assign io_oeb[9] = net235;
 assign io_out[18] = net45;
 assign io_out[19] = net46;
 assign io_out[1] = net42;
 assign io_out[20] = net47;
 assign io_out[21] = net48;
 assign io_out[22] = net49;
 assign io_out[23] = net50;
 assign io_out[24] = net51;
 assign io_out[25] = net52;
 assign io_out[26] = net53;
 assign io_out[27] = net54;
 assign io_out[28] = net55;
 assign io_out[29] = net56;
 assign io_out[2] = net43;
 assign io_out[30] = net57;
 assign io_out[31] = net58;
 assign io_out[32] = net59;
 assign io_out[33] = net60;
 assign io_out[34] = net61;
 assign io_out[35] = net62;
 assign io_out[36] = net63;
 assign io_out[37] = net64;
 assign io_out[3] = net44;
 assign la_data_out[0] = net65;
 assign la_data_out[100] = net133;
 assign la_data_out[101] = net134;
 assign la_data_out[102] = net135;
 assign la_data_out[103] = net136;
 assign la_data_out[104] = net137;
 assign la_data_out[105] = net138;
 assign la_data_out[106] = net139;
 assign la_data_out[107] = net140;
 assign la_data_out[108] = net141;
 assign la_data_out[109] = net142;
 assign la_data_out[10] = net75;
 assign la_data_out[110] = net143;
 assign la_data_out[111] = net144;
 assign la_data_out[112] = net145;
 assign la_data_out[113] = net146;
 assign la_data_out[114] = net147;
 assign la_data_out[115] = net148;
 assign la_data_out[116] = net149;
 assign la_data_out[117] = net150;
 assign la_data_out[118] = net151;
 assign la_data_out[119] = net152;
 assign la_data_out[11] = net76;
 assign la_data_out[120] = net153;
 assign la_data_out[121] = net154;
 assign la_data_out[122] = net155;
 assign la_data_out[123] = net156;
 assign la_data_out[124] = net157;
 assign la_data_out[125] = net158;
 assign la_data_out[126] = net159;
 assign la_data_out[127] = net160;
 assign la_data_out[12] = net77;
 assign la_data_out[13] = net78;
 assign la_data_out[14] = net79;
 assign la_data_out[15] = net80;
 assign la_data_out[16] = net81;
 assign la_data_out[17] = net82;
 assign la_data_out[18] = net83;
 assign la_data_out[19] = net84;
 assign la_data_out[1] = net66;
 assign la_data_out[20] = net85;
 assign la_data_out[21] = net86;
 assign la_data_out[22] = net87;
 assign la_data_out[23] = net88;
 assign la_data_out[24] = net89;
 assign la_data_out[25] = net90;
 assign la_data_out[26] = net91;
 assign la_data_out[27] = net92;
 assign la_data_out[28] = net93;
 assign la_data_out[29] = net94;
 assign la_data_out[2] = net67;
 assign la_data_out[30] = net95;
 assign la_data_out[31] = net96;
 assign la_data_out[3] = net68;
 assign la_data_out[4] = net69;
 assign la_data_out[5] = net70;
 assign la_data_out[64] = net97;
 assign la_data_out[65] = net98;
 assign la_data_out[66] = net99;
 assign la_data_out[67] = net100;
 assign la_data_out[68] = net101;
 assign la_data_out[69] = net102;
 assign la_data_out[6] = net71;
 assign la_data_out[70] = net103;
 assign la_data_out[71] = net104;
 assign la_data_out[72] = net105;
 assign la_data_out[73] = net106;
 assign la_data_out[74] = net107;
 assign la_data_out[75] = net108;
 assign la_data_out[76] = net109;
 assign la_data_out[77] = net110;
 assign la_data_out[78] = net111;
 assign la_data_out[79] = net112;
 assign la_data_out[7] = net72;
 assign la_data_out[80] = net113;
 assign la_data_out[81] = net114;
 assign la_data_out[82] = net115;
 assign la_data_out[83] = net116;
 assign la_data_out[84] = net117;
 assign la_data_out[85] = net118;
 assign la_data_out[86] = net119;
 assign la_data_out[87] = net120;
 assign la_data_out[88] = net121;
 assign la_data_out[89] = net122;
 assign la_data_out[8] = net73;
 assign la_data_out[90] = net123;
 assign la_data_out[91] = net124;
 assign la_data_out[92] = net125;
 assign la_data_out[93] = net126;
 assign la_data_out[94] = net127;
 assign la_data_out[95] = net128;
 assign la_data_out[96] = net129;
 assign la_data_out[97] = net130;
 assign la_data_out[98] = net131;
 assign la_data_out[99] = net132;
 assign la_data_out[9] = net74;
 assign wbs_ack_o = net161;
 assign wbs_dat_o[0] = net162;
 assign wbs_dat_o[10] = net172;
 assign wbs_dat_o[11] = net173;
 assign wbs_dat_o[12] = net174;
 assign wbs_dat_o[13] = net175;
 assign wbs_dat_o[14] = net176;
 assign wbs_dat_o[15] = net177;
 assign wbs_dat_o[16] = net178;
 assign wbs_dat_o[17] = net179;
 assign wbs_dat_o[18] = net180;
 assign wbs_dat_o[19] = net181;
 assign wbs_dat_o[1] = net163;
 assign wbs_dat_o[20] = net182;
 assign wbs_dat_o[21] = net183;
 assign wbs_dat_o[22] = net184;
 assign wbs_dat_o[23] = net185;
 assign wbs_dat_o[24] = net186;
 assign wbs_dat_o[25] = net187;
 assign wbs_dat_o[26] = net188;
 assign wbs_dat_o[27] = net189;
 assign wbs_dat_o[28] = net190;
 assign wbs_dat_o[29] = net191;
 assign wbs_dat_o[2] = net164;
 assign wbs_dat_o[30] = net192;
 assign wbs_dat_o[31] = net193;
 assign wbs_dat_o[3] = net165;
 assign wbs_dat_o[4] = net166;
 assign wbs_dat_o[5] = net167;
 assign wbs_dat_o[6] = net168;
 assign wbs_dat_o[7] = net169;
 assign wbs_dat_o[8] = net170;
 assign wbs_dat_o[9] = net171;
endmodule

