// This is the unpowered netlist.
module macro_15 (io_active,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input io_active;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net228;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net229;
 wire net257;
 wire net258;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net46;
 wire net47;
 wire net43;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net44;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net45;
 wire net66;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net76;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net77;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net67;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net68;
 wire net96;
 wire net97;
 wire net69;
 wire net70;
 wire net71;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net72;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net73;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net74;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net75;
 wire net162;
 wire net163;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net164;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net165;
 wire net193;
 wire net194;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;

 sky130_fd_sc_hd__inv_2 _157_ (.A(net1),
    .Y(_124_));
 sky130_fd_sc_hd__buf_4 _158_ (.A(net1),
    .X(_089_));
 sky130_fd_sc_hd__buf_4 _159_ (.A(_089_),
    .X(_090_));
 sky130_fd_sc_hd__inv_2 _160_ (.A(_090_),
    .Y(_123_));
 sky130_fd_sc_hd__inv_2 _161_ (.A(_090_),
    .Y(_122_));
 sky130_fd_sc_hd__inv_2 _162_ (.A(_090_),
    .Y(_121_));
 sky130_fd_sc_hd__inv_2 _163_ (.A(_090_),
    .Y(_120_));
 sky130_fd_sc_hd__inv_2 _164_ (.A(_090_),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _165_ (.A(_090_),
    .Y(_118_));
 sky130_fd_sc_hd__inv_2 _166_ (.A(_090_),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _167_ (.A(_090_),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _168_ (.A(_090_),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _169_ (.A(_090_),
    .Y(_114_));
 sky130_fd_sc_hd__buf_4 _170_ (.A(_089_),
    .X(_091_));
 sky130_fd_sc_hd__inv_2 _171_ (.A(_091_),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _172_ (.A(_091_),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _173_ (.A(_091_),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _174_ (.A(_091_),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _175_ (.A(_091_),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _176_ (.A(_091_),
    .Y(_108_));
 sky130_fd_sc_hd__inv_2 _177_ (.A(_091_),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _178_ (.A(_091_),
    .Y(_106_));
 sky130_fd_sc_hd__inv_2 _179_ (.A(_091_),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _180_ (.A(_091_),
    .Y(_104_));
 sky130_fd_sc_hd__buf_4 _181_ (.A(_089_),
    .X(_092_));
 sky130_fd_sc_hd__inv_2 _182_ (.A(_092_),
    .Y(_103_));
 sky130_fd_sc_hd__inv_2 _183_ (.A(_092_),
    .Y(_102_));
 sky130_fd_sc_hd__inv_2 _184_ (.A(_092_),
    .Y(_101_));
 sky130_fd_sc_hd__inv_2 _185_ (.A(_092_),
    .Y(_100_));
 sky130_fd_sc_hd__inv_2 _186_ (.A(_092_),
    .Y(_099_));
 sky130_fd_sc_hd__inv_2 _187_ (.A(_092_),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _188_ (.A(_092_),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _189_ (.A(_092_),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _190_ (.A(_092_),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _191_ (.A(_092_),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _192_ (.A(_089_),
    .Y(_093_));
 sky130_fd_sc_hd__nand2b_1 _193_ (.A_N(net19),
    .B(net18),
    .Y(_000_));
 sky130_fd_sc_hd__o31a_1 _194_ (.A1(net8),
    .A2(net6),
    .A3(net7),
    .B1(_000_),
    .X(_001_));
 sky130_fd_sc_hd__xnor2_1 _195_ (.A(net9),
    .B(_001_),
    .Y(_002_));
 sky130_fd_sc_hd__or2_1 _196_ (.A(net5),
    .B(_002_),
    .X(_003_));
 sky130_fd_sc_hd__o21a_1 _197_ (.A1(net6),
    .A2(net7),
    .B1(_000_),
    .X(_004_));
 sky130_fd_sc_hd__xnor2_1 _198_ (.A(net8),
    .B(_004_),
    .Y(_005_));
 sky130_fd_sc_hd__or2_1 _199_ (.A(net4),
    .B(_005_),
    .X(_006_));
 sky130_fd_sc_hd__nand3b_1 _200_ (.A_N(net7),
    .B(_000_),
    .C(net6),
    .Y(_007_));
 sky130_fd_sc_hd__a21bo_1 _201_ (.A1(net6),
    .A2(_000_),
    .B1_N(net7),
    .X(_008_));
 sky130_fd_sc_hd__a21o_1 _202_ (.A1(_007_),
    .A2(_008_),
    .B1(net3),
    .X(_009_));
 sky130_fd_sc_hd__or2b_1 _203_ (.A(net2),
    .B_N(net6),
    .X(_010_));
 sky130_fd_sc_hd__and3_1 _204_ (.A(net3),
    .B(_007_),
    .C(_008_),
    .X(_011_));
 sky130_fd_sc_hd__a21o_1 _205_ (.A1(_009_),
    .A2(_010_),
    .B1(_011_),
    .X(_012_));
 sky130_fd_sc_hd__and2_1 _206_ (.A(net5),
    .B(_002_),
    .X(_013_));
 sky130_fd_sc_hd__and2_1 _207_ (.A(net4),
    .B(_005_),
    .X(_014_));
 sky130_fd_sc_hd__a211o_1 _208_ (.A1(_006_),
    .A2(_012_),
    .B1(_013_),
    .C1(_014_),
    .X(_015_));
 sky130_fd_sc_hd__a21oi_1 _209_ (.A1(net9),
    .A2(_000_),
    .B1(_001_),
    .Y(_016_));
 sky130_fd_sc_hd__a21oi_1 _210_ (.A1(_003_),
    .A2(_015_),
    .B1(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__a31o_1 _211_ (.A1(_016_),
    .A2(_003_),
    .A3(_015_),
    .B1(net19),
    .X(_018_));
 sky130_fd_sc_hd__or2_1 _212_ (.A(_017_),
    .B(_018_),
    .X(_019_));
 sky130_fd_sc_hd__nand2b_1 _213_ (.A_N(net21),
    .B(net20),
    .Y(_020_));
 sky130_fd_sc_hd__o31a_1 _214_ (.A1(net16),
    .A2(net14),
    .A3(net15),
    .B1(_020_),
    .X(_021_));
 sky130_fd_sc_hd__xnor2_1 _215_ (.A(net17),
    .B(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__or2_1 _216_ (.A(net13),
    .B(_022_),
    .X(_023_));
 sky130_fd_sc_hd__o21a_1 _217_ (.A1(net14),
    .A2(net15),
    .B1(_020_),
    .X(_024_));
 sky130_fd_sc_hd__xnor2_1 _218_ (.A(net16),
    .B(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__or2_1 _219_ (.A(net12),
    .B(_025_),
    .X(_026_));
 sky130_fd_sc_hd__nand3b_1 _220_ (.A_N(net15),
    .B(_020_),
    .C(net14),
    .Y(_027_));
 sky130_fd_sc_hd__a21bo_1 _221_ (.A1(net14),
    .A2(_020_),
    .B1_N(net15),
    .X(_028_));
 sky130_fd_sc_hd__a21o_1 _222_ (.A1(_027_),
    .A2(_028_),
    .B1(net11),
    .X(_029_));
 sky130_fd_sc_hd__or2b_1 _223_ (.A(net10),
    .B_N(net14),
    .X(_030_));
 sky130_fd_sc_hd__and3_1 _224_ (.A(net11),
    .B(_027_),
    .C(_028_),
    .X(_031_));
 sky130_fd_sc_hd__a21o_1 _225_ (.A1(_029_),
    .A2(_030_),
    .B1(_031_),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _226_ (.A(net13),
    .B(_022_),
    .X(_033_));
 sky130_fd_sc_hd__and2_1 _227_ (.A(net12),
    .B(_025_),
    .X(_034_));
 sky130_fd_sc_hd__a211o_1 _228_ (.A1(_026_),
    .A2(_032_),
    .B1(_033_),
    .C1(_034_),
    .X(_035_));
 sky130_fd_sc_hd__a21oi_1 _229_ (.A1(net17),
    .A2(_020_),
    .B1(_021_),
    .Y(_036_));
 sky130_fd_sc_hd__a21oi_1 _230_ (.A1(_023_),
    .A2(_035_),
    .B1(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__a31o_1 _231_ (.A1(_036_),
    .A2(_023_),
    .A3(_035_),
    .B1(net21),
    .X(_038_));
 sky130_fd_sc_hd__or2_1 _232_ (.A(_037_),
    .B(_038_),
    .X(_039_));
 sky130_fd_sc_hd__nor3_2 _233_ (.A(_124_),
    .B(_037_),
    .C(_038_),
    .Y(net31));
 sky130_fd_sc_hd__nor3_1 _234_ (.A(_124_),
    .B(_017_),
    .C(_018_),
    .Y(net32));
 sky130_fd_sc_hd__o22a_1 _235_ (.A1(_019_),
    .A2(_039_),
    .B1(net31),
    .B2(net32),
    .X(net22));
 sky130_fd_sc_hd__inv_2 _236_ (.A(net19),
    .Y(_040_));
 sky130_fd_sc_hd__o2bb2a_1 _237_ (.A1_N(net6),
    .A2_N(net2),
    .B1(_040_),
    .B2(net18),
    .X(_041_));
 sky130_fd_sc_hd__o21a_1 _238_ (.A1(net6),
    .A2(net2),
    .B1(_041_),
    .X(_042_));
 sky130_fd_sc_hd__a31o_1 _239_ (.A1(net6),
    .A2(net19),
    .A3(net2),
    .B1(_042_),
    .X(_043_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(net21),
    .Y(_044_));
 sky130_fd_sc_hd__o2bb2a_1 _241_ (.A1_N(net14),
    .A2_N(net10),
    .B1(_044_),
    .B2(net20),
    .X(_045_));
 sky130_fd_sc_hd__o21a_1 _242_ (.A1(net14),
    .A2(net10),
    .B1(_045_),
    .X(_046_));
 sky130_fd_sc_hd__a31o_1 _243_ (.A1(net14),
    .A2(net21),
    .A3(net10),
    .B1(_046_),
    .X(_047_));
 sky130_fd_sc_hd__and2_1 _244_ (.A(_089_),
    .B(_047_),
    .X(_048_));
 sky130_fd_sc_hd__clkbuf_1 _245_ (.A(_048_),
    .X(net23));
 sky130_fd_sc_hd__and2_1 _246_ (.A(_089_),
    .B(_043_),
    .X(_049_));
 sky130_fd_sc_hd__clkbuf_1 _247_ (.A(_049_),
    .X(net27));
 sky130_fd_sc_hd__o2bb2a_1 _248_ (.A1_N(_043_),
    .A2_N(_047_),
    .B1(net23),
    .B2(net27),
    .X(net33));
 sky130_fd_sc_hd__or2b_1 _249_ (.A(_011_),
    .B_N(_009_),
    .X(_050_));
 sky130_fd_sc_hd__xnor2_1 _250_ (.A(_050_),
    .B(_010_),
    .Y(_051_));
 sky130_fd_sc_hd__o21a_1 _251_ (.A1(net7),
    .A2(net18),
    .B1(net3),
    .X(_052_));
 sky130_fd_sc_hd__a211o_1 _252_ (.A1(net7),
    .A2(net18),
    .B1(_040_),
    .C1(_052_),
    .X(_053_));
 sky130_fd_sc_hd__o21a_1 _253_ (.A1(net19),
    .A2(_051_),
    .B1(_053_),
    .X(_054_));
 sky130_fd_sc_hd__or2b_1 _254_ (.A(_031_),
    .B_N(_029_),
    .X(_055_));
 sky130_fd_sc_hd__xnor2_1 _255_ (.A(_055_),
    .B(_030_),
    .Y(_056_));
 sky130_fd_sc_hd__o21a_1 _256_ (.A1(net15),
    .A2(net20),
    .B1(net11),
    .X(_057_));
 sky130_fd_sc_hd__a211o_1 _257_ (.A1(net15),
    .A2(net20),
    .B1(_044_),
    .C1(_057_),
    .X(_058_));
 sky130_fd_sc_hd__o21a_1 _258_ (.A1(net21),
    .A2(_056_),
    .B1(_058_),
    .X(_059_));
 sky130_fd_sc_hd__and2_1 _259_ (.A(_089_),
    .B(_059_),
    .X(_060_));
 sky130_fd_sc_hd__clkbuf_1 _260_ (.A(_060_),
    .X(net24));
 sky130_fd_sc_hd__and2_1 _261_ (.A(_089_),
    .B(_054_),
    .X(_061_));
 sky130_fd_sc_hd__clkbuf_1 _262_ (.A(_061_),
    .X(net28));
 sky130_fd_sc_hd__o2bb2a_1 _263_ (.A1_N(_054_),
    .A2_N(_059_),
    .B1(net24),
    .B2(net28),
    .X(net34));
 sky130_fd_sc_hd__a21o_1 _264_ (.A1(net18),
    .A2(net4),
    .B1(net8),
    .X(_062_));
 sky130_fd_sc_hd__or2_1 _265_ (.A(net18),
    .B(net4),
    .X(_063_));
 sky130_fd_sc_hd__xor2_1 _266_ (.A(net4),
    .B(_005_),
    .X(_064_));
 sky130_fd_sc_hd__or2_1 _267_ (.A(_064_),
    .B(_012_),
    .X(_065_));
 sky130_fd_sc_hd__a21oi_1 _268_ (.A1(_064_),
    .A2(_012_),
    .B1(net19),
    .Y(_066_));
 sky130_fd_sc_hd__a32o_1 _269_ (.A1(net19),
    .A2(_062_),
    .A3(_063_),
    .B1(_065_),
    .B2(_066_),
    .X(_067_));
 sky130_fd_sc_hd__a21o_1 _270_ (.A1(net20),
    .A2(net12),
    .B1(net16),
    .X(_068_));
 sky130_fd_sc_hd__or2_1 _271_ (.A(net20),
    .B(net12),
    .X(_069_));
 sky130_fd_sc_hd__xor2_1 _272_ (.A(net12),
    .B(_025_),
    .X(_070_));
 sky130_fd_sc_hd__or2_1 _273_ (.A(_070_),
    .B(_032_),
    .X(_071_));
 sky130_fd_sc_hd__a21oi_1 _274_ (.A1(_070_),
    .A2(_032_),
    .B1(net21),
    .Y(_072_));
 sky130_fd_sc_hd__a32o_1 _275_ (.A1(net21),
    .A2(_068_),
    .A3(_069_),
    .B1(_071_),
    .B2(_072_),
    .X(_073_));
 sky130_fd_sc_hd__and2_1 _276_ (.A(net1),
    .B(_073_),
    .X(_074_));
 sky130_fd_sc_hd__clkbuf_1 _277_ (.A(_074_),
    .X(net25));
 sky130_fd_sc_hd__and2_1 _278_ (.A(_089_),
    .B(_067_),
    .X(_075_));
 sky130_fd_sc_hd__clkbuf_1 _279_ (.A(_075_),
    .X(net29));
 sky130_fd_sc_hd__o2bb2a_1 _280_ (.A1_N(_067_),
    .A2_N(_073_),
    .B1(net25),
    .B2(net29),
    .X(net35));
 sky130_fd_sc_hd__a21oi_1 _281_ (.A1(_006_),
    .A2(_012_),
    .B1(_014_),
    .Y(_076_));
 sky130_fd_sc_hd__and2b_1 _282_ (.A_N(_013_),
    .B(_003_),
    .X(_077_));
 sky130_fd_sc_hd__xnor2_1 _283_ (.A(_076_),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__nor2_1 _284_ (.A(net19),
    .B(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__o21a_1 _285_ (.A1(net9),
    .A2(net18),
    .B1(net5),
    .X(_080_));
 sky130_fd_sc_hd__a21o_1 _286_ (.A1(net9),
    .A2(net18),
    .B1(_040_),
    .X(_081_));
 sky130_fd_sc_hd__nor2_1 _287_ (.A(_080_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__a21o_1 _288_ (.A1(_026_),
    .A2(_032_),
    .B1(_034_),
    .X(_083_));
 sky130_fd_sc_hd__and2b_1 _289_ (.A_N(_033_),
    .B(_023_),
    .X(_084_));
 sky130_fd_sc_hd__xnor2_1 _290_ (.A(_083_),
    .B(_084_),
    .Y(_085_));
 sky130_fd_sc_hd__o21a_1 _291_ (.A1(net17),
    .A2(net20),
    .B1(net13),
    .X(_086_));
 sky130_fd_sc_hd__a211oi_2 _292_ (.A1(net17),
    .A2(net20),
    .B1(_044_),
    .C1(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__a21o_1 _293_ (.A1(_044_),
    .A2(_085_),
    .B1(_087_),
    .X(_088_));
 sky130_fd_sc_hd__a211oi_2 _294_ (.A1(_044_),
    .A2(_085_),
    .B1(_087_),
    .C1(_124_),
    .Y(net26));
 sky130_fd_sc_hd__o221a_1 _295_ (.A1(net19),
    .A2(_078_),
    .B1(_080_),
    .B2(_081_),
    .C1(_089_),
    .X(net30));
 sky130_fd_sc_hd__o32a_1 _296_ (.A1(_079_),
    .A2(_082_),
    .A3(_088_),
    .B1(net26),
    .B2(net30),
    .X(net36));
 sky130_fd_sc_hd__conb_1 macro_15_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 macro_15_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 macro_15_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 macro_15_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 macro_15_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 macro_15_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 macro_15_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 macro_15_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 macro_15_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 macro_15_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 macro_15_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 macro_15_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 macro_15_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 macro_15_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 macro_15_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 macro_15_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 macro_15_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 macro_15_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 macro_15_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 macro_15_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 macro_15_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 macro_15_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 macro_15_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 macro_15_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 macro_15_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 macro_15_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 macro_15_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 macro_15_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 macro_15_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 macro_15_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 macro_15_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 macro_15_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 macro_15_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 macro_15_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 macro_15_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 macro_15_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 macro_15_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 macro_15_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 macro_15_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 macro_15_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 macro_15_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 macro_15_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 macro_15_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 macro_15_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 macro_15_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 macro_15_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 macro_15_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 macro_15_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 macro_15_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 macro_15_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 macro_15_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 macro_15_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 macro_15_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 macro_15_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 macro_15_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 macro_15_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 macro_15_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 macro_15_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 macro_15_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 macro_15_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 macro_15_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 macro_15_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 macro_15_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 macro_15_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 macro_15_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 macro_15_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 macro_15_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 macro_15_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 macro_15_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 macro_15_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 macro_15_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 macro_15_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 macro_15_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 macro_15_111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 macro_15_112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 macro_15_113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 macro_15_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 macro_15_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 macro_15_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 macro_15_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 macro_15_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 macro_15_119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 macro_15_120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 macro_15_121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 macro_15_122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 macro_15_123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 macro_15_124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 macro_15_125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 macro_15_126 (.LO(net126));
 sky130_fd_sc_hd__conb_1 macro_15_127 (.LO(net127));
 sky130_fd_sc_hd__conb_1 macro_15_128 (.LO(net128));
 sky130_fd_sc_hd__conb_1 macro_15_129 (.LO(net129));
 sky130_fd_sc_hd__conb_1 macro_15_130 (.LO(net130));
 sky130_fd_sc_hd__conb_1 macro_15_131 (.LO(net131));
 sky130_fd_sc_hd__conb_1 macro_15_132 (.LO(net132));
 sky130_fd_sc_hd__conb_1 macro_15_133 (.LO(net133));
 sky130_fd_sc_hd__conb_1 macro_15_134 (.LO(net134));
 sky130_fd_sc_hd__conb_1 macro_15_135 (.LO(net135));
 sky130_fd_sc_hd__conb_1 macro_15_136 (.LO(net136));
 sky130_fd_sc_hd__conb_1 macro_15_137 (.LO(net137));
 sky130_fd_sc_hd__conb_1 macro_15_138 (.LO(net138));
 sky130_fd_sc_hd__conb_1 macro_15_139 (.LO(net139));
 sky130_fd_sc_hd__conb_1 macro_15_140 (.LO(net140));
 sky130_fd_sc_hd__conb_1 macro_15_141 (.LO(net141));
 sky130_fd_sc_hd__conb_1 macro_15_142 (.LO(net142));
 sky130_fd_sc_hd__conb_1 macro_15_143 (.LO(net143));
 sky130_fd_sc_hd__conb_1 macro_15_144 (.LO(net144));
 sky130_fd_sc_hd__conb_1 macro_15_145 (.LO(net145));
 sky130_fd_sc_hd__conb_1 macro_15_146 (.LO(net146));
 sky130_fd_sc_hd__conb_1 macro_15_147 (.LO(net147));
 sky130_fd_sc_hd__conb_1 macro_15_148 (.LO(net148));
 sky130_fd_sc_hd__conb_1 macro_15_149 (.LO(net149));
 sky130_fd_sc_hd__conb_1 macro_15_150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 macro_15_151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 macro_15_152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 macro_15_153 (.LO(net153));
 sky130_fd_sc_hd__conb_1 macro_15_154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 macro_15_155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 macro_15_156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 macro_15_157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 macro_15_158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 macro_15_159 (.LO(net159));
 sky130_fd_sc_hd__conb_1 macro_15_160 (.LO(net160));
 sky130_fd_sc_hd__conb_1 macro_15_161 (.LO(net161));
 sky130_fd_sc_hd__conb_1 macro_15_162 (.LO(net162));
 sky130_fd_sc_hd__conb_1 macro_15_163 (.LO(net163));
 sky130_fd_sc_hd__conb_1 macro_15_164 (.LO(net164));
 sky130_fd_sc_hd__conb_1 macro_15_165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 macro_15_166 (.LO(net166));
 sky130_fd_sc_hd__conb_1 macro_15_167 (.LO(net167));
 sky130_fd_sc_hd__conb_1 macro_15_168 (.LO(net168));
 sky130_fd_sc_hd__conb_1 macro_15_169 (.LO(net169));
 sky130_fd_sc_hd__conb_1 macro_15_170 (.LO(net170));
 sky130_fd_sc_hd__conb_1 macro_15_171 (.LO(net171));
 sky130_fd_sc_hd__conb_1 macro_15_172 (.LO(net172));
 sky130_fd_sc_hd__conb_1 macro_15_173 (.LO(net173));
 sky130_fd_sc_hd__conb_1 macro_15_174 (.LO(net174));
 sky130_fd_sc_hd__conb_1 macro_15_175 (.LO(net175));
 sky130_fd_sc_hd__conb_1 macro_15_176 (.LO(net176));
 sky130_fd_sc_hd__conb_1 macro_15_177 (.LO(net177));
 sky130_fd_sc_hd__conb_1 macro_15_178 (.LO(net178));
 sky130_fd_sc_hd__conb_1 macro_15_179 (.LO(net179));
 sky130_fd_sc_hd__conb_1 macro_15_180 (.LO(net180));
 sky130_fd_sc_hd__conb_1 macro_15_181 (.LO(net181));
 sky130_fd_sc_hd__conb_1 macro_15_182 (.LO(net182));
 sky130_fd_sc_hd__conb_1 macro_15_183 (.LO(net183));
 sky130_fd_sc_hd__conb_1 macro_15_184 (.LO(net184));
 sky130_fd_sc_hd__conb_1 macro_15_185 (.LO(net185));
 sky130_fd_sc_hd__conb_1 macro_15_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 macro_15_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 macro_15_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 macro_15_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 macro_15_190 (.LO(net190));
 sky130_fd_sc_hd__conb_1 macro_15_191 (.LO(net191));
 sky130_fd_sc_hd__conb_1 macro_15_192 (.LO(net192));
 sky130_fd_sc_hd__conb_1 macro_15_193 (.LO(net193));
 sky130_fd_sc_hd__conb_1 _519__194 (.LO(net194));
 sky130_fd_sc_hd__conb_1 _520__195 (.LO(net195));
 sky130_fd_sc_hd__conb_1 _521__196 (.LO(net196));
 sky130_fd_sc_hd__conb_1 _522__197 (.LO(net197));
 sky130_fd_sc_hd__conb_1 _523__198 (.LO(net198));
 sky130_fd_sc_hd__conb_1 _524__199 (.LO(net199));
 sky130_fd_sc_hd__conb_1 _525__200 (.LO(net200));
 sky130_fd_sc_hd__conb_1 _526__201 (.LO(net201));
 sky130_fd_sc_hd__conb_1 _527__202 (.LO(net202));
 sky130_fd_sc_hd__conb_1 _528__203 (.LO(net203));
 sky130_fd_sc_hd__conb_1 _529__204 (.LO(net204));
 sky130_fd_sc_hd__conb_1 _530__205 (.LO(net205));
 sky130_fd_sc_hd__conb_1 _531__206 (.LO(net206));
 sky130_fd_sc_hd__conb_1 _532__207 (.LO(net207));
 sky130_fd_sc_hd__conb_1 _533__208 (.LO(net208));
 sky130_fd_sc_hd__conb_1 _534__209 (.LO(net209));
 sky130_fd_sc_hd__conb_1 _535__210 (.LO(net210));
 sky130_fd_sc_hd__conb_1 _536__211 (.LO(net211));
 sky130_fd_sc_hd__conb_1 _537__212 (.LO(net212));
 sky130_fd_sc_hd__conb_1 _538__213 (.LO(net213));
 sky130_fd_sc_hd__conb_1 _539__214 (.LO(net214));
 sky130_fd_sc_hd__conb_1 _540__215 (.LO(net215));
 sky130_fd_sc_hd__conb_1 _541__216 (.LO(net216));
 sky130_fd_sc_hd__conb_1 _542__217 (.LO(net217));
 sky130_fd_sc_hd__conb_1 _543__218 (.LO(net218));
 sky130_fd_sc_hd__conb_1 _544__219 (.LO(net219));
 sky130_fd_sc_hd__conb_1 _545__220 (.LO(net220));
 sky130_fd_sc_hd__conb_1 _546__221 (.LO(net221));
 sky130_fd_sc_hd__conb_1 _547__222 (.LO(net222));
 sky130_fd_sc_hd__conb_1 _548__223 (.LO(net223));
 sky130_fd_sc_hd__conb_1 _549__224 (.LO(net224));
 sky130_fd_sc_hd__conb_1 _550__225 (.LO(net225));
 sky130_fd_sc_hd__conb_1 macro_15_226 (.LO(net226));
 sky130_fd_sc_hd__conb_1 macro_15_227 (.LO(net227));
 sky130_fd_sc_hd__conb_1 macro_15_228 (.LO(net228));
 sky130_fd_sc_hd__conb_1 macro_15_229 (.LO(net229));
 sky130_fd_sc_hd__conb_1 macro_15_230 (.LO(net230));
 sky130_fd_sc_hd__conb_1 macro_15_231 (.LO(net231));
 sky130_fd_sc_hd__conb_1 macro_15_232 (.LO(net232));
 sky130_fd_sc_hd__conb_1 macro_15_233 (.LO(net233));
 sky130_fd_sc_hd__conb_1 macro_15_234 (.LO(net234));
 sky130_fd_sc_hd__conb_1 macro_15_235 (.LO(net235));
 sky130_fd_sc_hd__conb_1 macro_15_236 (.LO(net236));
 sky130_fd_sc_hd__conb_1 macro_15_237 (.LO(net237));
 sky130_fd_sc_hd__conb_1 macro_15_238 (.LO(net238));
 sky130_fd_sc_hd__conb_1 macro_15_239 (.LO(net239));
 sky130_fd_sc_hd__conb_1 macro_15_240 (.LO(net240));
 sky130_fd_sc_hd__conb_1 macro_15_241 (.LO(net241));
 sky130_fd_sc_hd__conb_1 macro_15_242 (.LO(net242));
 sky130_fd_sc_hd__conb_1 macro_15_243 (.LO(net243));
 sky130_fd_sc_hd__conb_1 macro_15_244 (.LO(net244));
 sky130_fd_sc_hd__conb_1 macro_15_245 (.LO(net245));
 sky130_fd_sc_hd__conb_1 macro_15_246 (.LO(net246));
 sky130_fd_sc_hd__conb_1 macro_15_247 (.LO(net247));
 sky130_fd_sc_hd__conb_1 macro_15_248 (.LO(net248));
 sky130_fd_sc_hd__conb_1 macro_15_249 (.LO(net249));
 sky130_fd_sc_hd__conb_1 macro_15_250 (.LO(net250));
 sky130_fd_sc_hd__conb_1 macro_15_251 (.LO(net251));
 sky130_fd_sc_hd__conb_1 macro_15_252 (.LO(net252));
 sky130_fd_sc_hd__conb_1 macro_15_253 (.LO(net253));
 sky130_fd_sc_hd__conb_1 macro_15_254 (.LO(net254));
 sky130_fd_sc_hd__conb_1 macro_15_255 (.LO(net255));
 sky130_fd_sc_hd__conb_1 macro_15_256 (.LO(net256));
 sky130_fd_sc_hd__conb_1 macro_15_257 (.LO(net257));
 sky130_fd_sc_hd__conb_1 macro_15_258 (.LO(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__C1 (.DIODE(_089_));
 sky130_fd_sc_hd__ebufn_8 _519_ (.A(net194),
    .TE_B(_093_),
    .Z(la_data_out[32]));
 sky130_fd_sc_hd__ebufn_8 _520_ (.A(net195),
    .TE_B(_094_),
    .Z(la_data_out[33]));
 sky130_fd_sc_hd__ebufn_8 _521_ (.A(net196),
    .TE_B(_095_),
    .Z(la_data_out[34]));
 sky130_fd_sc_hd__ebufn_8 _522_ (.A(net197),
    .TE_B(_096_),
    .Z(la_data_out[35]));
 sky130_fd_sc_hd__ebufn_8 _523_ (.A(net198),
    .TE_B(_097_),
    .Z(la_data_out[36]));
 sky130_fd_sc_hd__ebufn_8 _524_ (.A(net199),
    .TE_B(_098_),
    .Z(la_data_out[37]));
 sky130_fd_sc_hd__ebufn_8 _525_ (.A(net200),
    .TE_B(_099_),
    .Z(la_data_out[38]));
 sky130_fd_sc_hd__ebufn_8 _526_ (.A(net201),
    .TE_B(_100_),
    .Z(la_data_out[39]));
 sky130_fd_sc_hd__ebufn_8 _527_ (.A(net202),
    .TE_B(_101_),
    .Z(la_data_out[40]));
 sky130_fd_sc_hd__ebufn_8 _528_ (.A(net203),
    .TE_B(_102_),
    .Z(la_data_out[41]));
 sky130_fd_sc_hd__ebufn_8 _529_ (.A(net204),
    .TE_B(_103_),
    .Z(la_data_out[42]));
 sky130_fd_sc_hd__ebufn_8 _530_ (.A(net205),
    .TE_B(_104_),
    .Z(la_data_out[43]));
 sky130_fd_sc_hd__ebufn_8 _531_ (.A(net206),
    .TE_B(_105_),
    .Z(la_data_out[44]));
 sky130_fd_sc_hd__ebufn_8 _532_ (.A(net207),
    .TE_B(_106_),
    .Z(la_data_out[45]));
 sky130_fd_sc_hd__ebufn_8 _533_ (.A(net208),
    .TE_B(_107_),
    .Z(la_data_out[46]));
 sky130_fd_sc_hd__ebufn_8 _534_ (.A(net209),
    .TE_B(_108_),
    .Z(la_data_out[47]));
 sky130_fd_sc_hd__ebufn_8 _535_ (.A(net210),
    .TE_B(_109_),
    .Z(la_data_out[48]));
 sky130_fd_sc_hd__ebufn_8 _536_ (.A(net211),
    .TE_B(_110_),
    .Z(la_data_out[49]));
 sky130_fd_sc_hd__ebufn_8 _537_ (.A(net212),
    .TE_B(_111_),
    .Z(la_data_out[50]));
 sky130_fd_sc_hd__ebufn_8 _538_ (.A(net213),
    .TE_B(_112_),
    .Z(la_data_out[51]));
 sky130_fd_sc_hd__ebufn_8 _539_ (.A(net214),
    .TE_B(_113_),
    .Z(la_data_out[52]));
 sky130_fd_sc_hd__ebufn_8 _540_ (.A(net215),
    .TE_B(_114_),
    .Z(la_data_out[53]));
 sky130_fd_sc_hd__ebufn_8 _541_ (.A(net216),
    .TE_B(_115_),
    .Z(la_data_out[54]));
 sky130_fd_sc_hd__ebufn_8 _542_ (.A(net217),
    .TE_B(_116_),
    .Z(la_data_out[55]));
 sky130_fd_sc_hd__ebufn_8 _543_ (.A(net218),
    .TE_B(_117_),
    .Z(la_data_out[56]));
 sky130_fd_sc_hd__ebufn_8 _544_ (.A(net219),
    .TE_B(_118_),
    .Z(la_data_out[57]));
 sky130_fd_sc_hd__ebufn_8 _545_ (.A(net220),
    .TE_B(_119_),
    .Z(la_data_out[58]));
 sky130_fd_sc_hd__ebufn_8 _546_ (.A(net221),
    .TE_B(_120_),
    .Z(la_data_out[59]));
 sky130_fd_sc_hd__ebufn_8 _547_ (.A(net222),
    .TE_B(_121_),
    .Z(la_data_out[60]));
 sky130_fd_sc_hd__ebufn_8 _548_ (.A(net223),
    .TE_B(_122_),
    .Z(la_data_out[61]));
 sky130_fd_sc_hd__ebufn_8 _549_ (.A(net224),
    .TE_B(_123_),
    .Z(la_data_out[62]));
 sky130_fd_sc_hd__ebufn_8 _550_ (.A(net225),
    .TE_B(_124_),
    .Z(la_data_out[63]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_active),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[18]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[19]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(io_in[20]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[21]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[22]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(io_in[23]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(io_in[24]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(io_in[25]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(io_in[26]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(io_in[27]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(io_in[28]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(io_in[29]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(io_in[30]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(io_in[31]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(io_in[32]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(io_in[33]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(io_in[34]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(io_in[35]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(io_in[36]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(io_in[37]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(io_out[9]));
 sky130_fd_sc_hd__conb_1 macro_15_37 (.LO(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__278__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__261__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__259__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__246__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__170__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__159__A (.DIODE(_089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_active));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(io_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(io_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(io_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__157__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__286__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__285__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__265__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__284__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__269__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__253__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__236__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__A_N (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__274__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__231__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__A_N (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__B1 (.DIODE(net31));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_621 ();
 assign io_oeb[0] = net226;
 assign io_oeb[10] = net236;
 assign io_oeb[11] = net237;
 assign io_oeb[12] = net238;
 assign io_oeb[13] = net239;
 assign io_oeb[14] = net240;
 assign io_oeb[15] = net241;
 assign io_oeb[16] = net242;
 assign io_oeb[17] = net243;
 assign io_oeb[18] = net244;
 assign io_oeb[19] = net245;
 assign io_oeb[1] = net227;
 assign io_oeb[20] = net246;
 assign io_oeb[21] = net247;
 assign io_oeb[22] = net248;
 assign io_oeb[23] = net249;
 assign io_oeb[24] = net250;
 assign io_oeb[25] = net251;
 assign io_oeb[26] = net252;
 assign io_oeb[27] = net253;
 assign io_oeb[28] = net254;
 assign io_oeb[29] = net255;
 assign io_oeb[2] = net228;
 assign io_oeb[30] = net256;
 assign io_oeb[31] = net257;
 assign io_oeb[32] = net258;
 assign io_oeb[33] = net37;
 assign io_oeb[34] = net38;
 assign io_oeb[35] = net39;
 assign io_oeb[36] = net40;
 assign io_oeb[37] = net41;
 assign io_oeb[3] = net229;
 assign io_oeb[4] = net230;
 assign io_oeb[5] = net231;
 assign io_oeb[6] = net232;
 assign io_oeb[7] = net233;
 assign io_oeb[8] = net234;
 assign io_oeb[9] = net235;
 assign io_out[18] = net45;
 assign io_out[19] = net46;
 assign io_out[1] = net42;
 assign io_out[20] = net47;
 assign io_out[21] = net48;
 assign io_out[22] = net49;
 assign io_out[23] = net50;
 assign io_out[24] = net51;
 assign io_out[25] = net52;
 assign io_out[26] = net53;
 assign io_out[27] = net54;
 assign io_out[28] = net55;
 assign io_out[29] = net56;
 assign io_out[2] = net43;
 assign io_out[30] = net57;
 assign io_out[31] = net58;
 assign io_out[32] = net59;
 assign io_out[33] = net60;
 assign io_out[34] = net61;
 assign io_out[35] = net62;
 assign io_out[36] = net63;
 assign io_out[37] = net64;
 assign io_out[3] = net44;
 assign la_data_out[0] = net65;
 assign la_data_out[100] = net133;
 assign la_data_out[101] = net134;
 assign la_data_out[102] = net135;
 assign la_data_out[103] = net136;
 assign la_data_out[104] = net137;
 assign la_data_out[105] = net138;
 assign la_data_out[106] = net139;
 assign la_data_out[107] = net140;
 assign la_data_out[108] = net141;
 assign la_data_out[109] = net142;
 assign la_data_out[10] = net75;
 assign la_data_out[110] = net143;
 assign la_data_out[111] = net144;
 assign la_data_out[112] = net145;
 assign la_data_out[113] = net146;
 assign la_data_out[114] = net147;
 assign la_data_out[115] = net148;
 assign la_data_out[116] = net149;
 assign la_data_out[117] = net150;
 assign la_data_out[118] = net151;
 assign la_data_out[119] = net152;
 assign la_data_out[11] = net76;
 assign la_data_out[120] = net153;
 assign la_data_out[121] = net154;
 assign la_data_out[122] = net155;
 assign la_data_out[123] = net156;
 assign la_data_out[124] = net157;
 assign la_data_out[125] = net158;
 assign la_data_out[126] = net159;
 assign la_data_out[127] = net160;
 assign la_data_out[12] = net77;
 assign la_data_out[13] = net78;
 assign la_data_out[14] = net79;
 assign la_data_out[15] = net80;
 assign la_data_out[16] = net81;
 assign la_data_out[17] = net82;
 assign la_data_out[18] = net83;
 assign la_data_out[19] = net84;
 assign la_data_out[1] = net66;
 assign la_data_out[20] = net85;
 assign la_data_out[21] = net86;
 assign la_data_out[22] = net87;
 assign la_data_out[23] = net88;
 assign la_data_out[24] = net89;
 assign la_data_out[25] = net90;
 assign la_data_out[26] = net91;
 assign la_data_out[27] = net92;
 assign la_data_out[28] = net93;
 assign la_data_out[29] = net94;
 assign la_data_out[2] = net67;
 assign la_data_out[30] = net95;
 assign la_data_out[31] = net96;
 assign la_data_out[3] = net68;
 assign la_data_out[4] = net69;
 assign la_data_out[5] = net70;
 assign la_data_out[64] = net97;
 assign la_data_out[65] = net98;
 assign la_data_out[66] = net99;
 assign la_data_out[67] = net100;
 assign la_data_out[68] = net101;
 assign la_data_out[69] = net102;
 assign la_data_out[6] = net71;
 assign la_data_out[70] = net103;
 assign la_data_out[71] = net104;
 assign la_data_out[72] = net105;
 assign la_data_out[73] = net106;
 assign la_data_out[74] = net107;
 assign la_data_out[75] = net108;
 assign la_data_out[76] = net109;
 assign la_data_out[77] = net110;
 assign la_data_out[78] = net111;
 assign la_data_out[79] = net112;
 assign la_data_out[7] = net72;
 assign la_data_out[80] = net113;
 assign la_data_out[81] = net114;
 assign la_data_out[82] = net115;
 assign la_data_out[83] = net116;
 assign la_data_out[84] = net117;
 assign la_data_out[85] = net118;
 assign la_data_out[86] = net119;
 assign la_data_out[87] = net120;
 assign la_data_out[88] = net121;
 assign la_data_out[89] = net122;
 assign la_data_out[8] = net73;
 assign la_data_out[90] = net123;
 assign la_data_out[91] = net124;
 assign la_data_out[92] = net125;
 assign la_data_out[93] = net126;
 assign la_data_out[94] = net127;
 assign la_data_out[95] = net128;
 assign la_data_out[96] = net129;
 assign la_data_out[97] = net130;
 assign la_data_out[98] = net131;
 assign la_data_out[99] = net132;
 assign la_data_out[9] = net74;
 assign wbs_ack_o = net161;
 assign wbs_dat_o[0] = net162;
 assign wbs_dat_o[10] = net172;
 assign wbs_dat_o[11] = net173;
 assign wbs_dat_o[12] = net174;
 assign wbs_dat_o[13] = net175;
 assign wbs_dat_o[14] = net176;
 assign wbs_dat_o[15] = net177;
 assign wbs_dat_o[16] = net178;
 assign wbs_dat_o[17] = net179;
 assign wbs_dat_o[18] = net180;
 assign wbs_dat_o[19] = net181;
 assign wbs_dat_o[1] = net163;
 assign wbs_dat_o[20] = net182;
 assign wbs_dat_o[21] = net183;
 assign wbs_dat_o[22] = net184;
 assign wbs_dat_o[23] = net185;
 assign wbs_dat_o[24] = net186;
 assign wbs_dat_o[25] = net187;
 assign wbs_dat_o[26] = net188;
 assign wbs_dat_o[27] = net189;
 assign wbs_dat_o[28] = net190;
 assign wbs_dat_o[29] = net191;
 assign wbs_dat_o[2] = net164;
 assign wbs_dat_o[30] = net192;
 assign wbs_dat_o[31] = net193;
 assign wbs_dat_o[3] = net165;
 assign wbs_dat_o[4] = net166;
 assign wbs_dat_o[5] = net167;
 assign wbs_dat_o[6] = net168;
 assign wbs_dat_o[7] = net169;
 assign wbs_dat_o[8] = net170;
 assign wbs_dat_o[9] = net171;
endmodule

